��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<��������T�]NA��M �\���(�	Bu� �k�A�=���:����V5p�N�=J��s�U#(�W�Iޖ�2�0���d��&����V�3@�&�E ݊O�J�O:0l)W��:@�]*}-�i��P0�3�׀�����8�7:�����=Bjњt�p�0hC}�#ǯ�G{�.�P�ƨ�o<�?/?�N�n�*��i���,8q���+���_�o��˔:Q)�p���o���Ap=��+�_]�A>i�4��-b������S��z����uQ����s �N � �ʿ�f鷍f˼�XdL��O��lB�'���-Q����t4�Vݽc1�Z���d�����y�@��༱I� "
Us�t��	���0�
��;�]>�E�,̼�u҈;M����^O#�f�ʮ���mf�rb6����������>�8B�	X6�Fo#�j7.J W�/���
�2)��YO��}8H'��b~��b/'$���p�ʬ%�6�l�x^�ȳXl�9����f��iX��~��tS�@]I�Y {y��FSV��`�_���B��tZ_�|�n�#
�:�Ֆ�8�g���F���]m%�<�'3zc6s}E]t�����ѧH��J���QEŧڅ���Y���%�:��x#r����?dד��Runy�q!?�ɐ�;��&.��x�L?IhG�Q�fna�&��f}�Z��4�zq��Z����Y���#�ļ�4��u��6�uF*(Q�%8�㟆f�f*��H�&�>�D���CBF{���-�C��p+s�~ݞ����y@A:�:kB�N�bR�Ig���ѕ&�:I�(�iG�>o0b�(�,$uT{+����(��Nvo�E�@�/QJ�Ɓ��*p
���C�8��^���E��G^�}�����6�� I$�W�̗{�k"�M�c�k�@Q7�n`e�cds���˅G �y%�	/2��� /�:���n�V��Z��-�Hv���6^U�dvw*�*f`Cս�g�Ɗ���c��\�J[�4�Pӥ'��з���x����RTn�pr����Ǚ��闿Bj��>7)cwE�6J���Q��v��f�q-I&l�%I�G�!�ޟ&���H��F՛(�������j<DB<7w��u�,+?ϭ�}ad��u ��3�b3�d���b/8M��0�j$�/�G!E��[T�C=��Ь��U5��-���}ϖ�{Ƥ��z%]2q�os����!�*�c�y�Q���먺����H󋩥���*Y���A��E*�uD�Ȳ�]"��-6%�L� ~ �j�>�|�I���3�f ��|�^X��x��3�OJ�ʨ�c
&���_bC�G�Ip�\l���8ϡ��!�_�5U��X��Q�?e���zsLO��]�5)?P-�2�i��[��p��U���b[ �_�u��t�^�m2N�B?�r�C��i�1<^Ե���r��t=��%Z�(�%��$�^Yx��IT.$_�����P(.�vSs����(:Qԝ�f�:Ku9e�Z��<�o����%���%�N$?����[:�<B�s��{/���!b3��%Z�I�A�-����T������Hh�`�����F9�2"m�"0�!Z���Vߑ������������h狿���3ڙ�R/A�0�m�r�T.�y���ﾶڇ���A27�َT͈Ǝ�ڇ��u2@��̮�X�3!!�ѐ�/dT0EJ�� ���� 4���J
<�N_�H���,�k��J7�?��B�����[��2Hڈ��Ƿ�Ài%�9�pL��c�ϧ�Aj�h.�(I�P�'�_����A���~�?^�d�4�{uؖ��v��<	Y��Ϫ�.o(]<db�>��@�q�<]���J�
�����-�y�U9�}�&��a B���J��|�(����8N�?��6V�Jqɭq��	 w�= ��_ӝq%G-M�=�)x�����A��|7�%_�\�����3���@藳W�E�Q��,�d燴٢c	��	�����/(	}fh������ͻ��6B����܇v��`0����y�t���\E�`�LhHOT�*~ς~�=�l�˲�-�VD�5y��݅�'1�5��|�OC�*���⪥s��Q�̻]S���&Z�c��`���$)6oF�9ro�����bٺ��m
J�\�xTo�C+H�9�����d4��]<�b���"������՘{����]��l�J6=�<_���H���z�cq-m�����9߂y#��yz���>�s�QY�_��.��|[Lʧz��,�ƻeT�e������g��c)#��-�y�S�e�����:�p?�D=xz3����
<w|Qt'	dI�p�� ��wZ�P�r;װ�c���w���c(Bͣwӽ�tƚ�}�� ���FC����������M�G�Ć�i���D.+v���A{�óq�ҧX�4���pa�Ki���L��#}b�*WB��.����n�X��S�����[����$U��H�VG�Gq��]M�#�97w�"�ވ#Y2�/E؅��>��o��%m�3 3��,L[}�l��@�ާ�:���S�����F����H��:�[2���Z.e��T3���0�����Fe�u�X��hۜ�B��#馧~���j�>��e
Ǉ�N��p��C��N' �C�;�%_�v�.��Zt�����y#�;�ph4-�� P���=��X���T��N����nV඗蠁�3�a��\(�oP�F����
/��`��w3��M��Ѷ�c�3ϣE��_Z���T�t��ۤ�i��6&
���&GY�����Yar�3yA$�ԏc�k���<����F��#3`Ǫ���B.�t��!͡}���)`69�H�K����K2w�D�!ZPDd0�
���<��do�tmjȆ����m�E�4˛�:9�����3#4Y�[xfnm<�����B<ٙ����R��eq����L�k��:X*4̞�'K6�M��~�C�5���ߕejDF�V�k��BT[�)���1��nf8	�*7/ؾE���97nE����u ���Z�y�/kR?@�%u:����9s�l]��Y?�/V/[N��&@�w��4�j��#��{{���Q�B�v��n.�H��e�T��n ��4��k$Ta�>���?�"��ޠ��b|��~V}Z�%"�z���M��#�I[�!��P�4��\��#v�9m�ډ���R2���$%��[���'@���@}V�#�������22l[`q�2(;���&v��"����|���F��(��k���@+�`�����ϸl�w�GВ�?c�Lѻ����-+M~㌩�lWx�S�*�%��D����L�%