��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<������::A���� �\�7�ݡ�y׵��G^.R��C\K�xef1�SDs����G2�km�����I��
�[��-��3�oX�by[���_K,�����J.ċS-���Q`�oS��{�������2���A�,N�`�n��e��>���b�EԞ�x�_��)D]�H��H�c)���#B(9�������ʒ�AQ����(l<�P@1Nmi+�W� 4%�0������޿��z�;�uU���C�ܴ�ѓ̱�y�Qx������d����f:w���4�������k!��Vx�(����+ʑ~�,.\Eޥmq$�ۄ�OQg��S��,�,�6ǘ�n����J:�]Y�>���8h��]K�"F��;�Ѐ�
��ml���+mZo8��E`�U��UIVN%�5�u�� ����<�����蟧L��b�WyɊϛ 
���.�u�ࢯ�����/k�4L��s����%�p�,g�����yg����w������3���;�'I����ŰKڒ�`l�Fu?Y���Bh+�w����D�r���F?���l���=P���a�XS�:�^��/��m�~��Y�Z�LP?cM�JZٗ�S˚���1-�]��H�Ni��(}��ьg��N��EG�p��/**�����0�2uu�����w���1���!���ª�+%�g}FZ5� �����֡>]W�:�6	��2qߜ �T����-����L
,�Q��K���E��ԁ��H�
�B��F=����}Uht��	!�5,�u�X(�*�6���������պ�iDKn�b���;��C�����=�l>8
�wm�M$��΃�솶}%������̷|��OU�V;vV��2ۣ���I7����S0P��`�܊����(�J��|�J*�۟hj��X,�4�gC����uZ���q�A�	�R�Q�[�����>ő��ǿ�� ?����]�AK[�78���}s�Ƭ����X�w ����q���oV�x1p�;��o��R����X6�=���<��U�P7�Ψ��"'R={�|7~�N�ΒIHz%�@��W6o�����%H��1܊�����^)=d	�N�8�A���y��^���%e������U��uy��o7I	J������"�������T���u���_V�67�ȭ�?i�D��
��&W���X�)�n����N̚�ݧ�6W���o.�ݹ7�� |3��j�T�X�/r7	Ƿ����6��]�� ��y�iL2	�Ge�C�E{h�L��)�X�f����5��	��k\<=b�/v�L�5�
#h����l��.I����n�H:�?�EȞ䠾��j�i�6����,B�N�����j���0D��tZ]X�w
�@Q�O���F5
#��+�nz:��zD��ՙ����%���8���"��#zOwmzivu��i�u7Bi��6P�wH�*��X_9 /u+>p
������p�3�e9�%�p��/pF�U6�q��R�kc�kvJ�f���ޤ{ɔ�G��$��@�Ɏ,�VSx��al�e����=�����͵^�n#��vM�_��P��8������o�R�;�OP'է2�oh�g�qgHvCh�Ҩo*7��ċ�S}���̌�@���5�(i!7���5Cr�QzcN����e2ʻ��\a��1�܋�O�t����������y��!�Ԕ�}q�A�5҃x��g���ɢ�a���4�8����S�s�`�a��I���DZ�ȕ�z��.���G�:a_h]̸����h�kM��_e=��=ͯ��s�s���Ț��6�y�$]��LL�^�Yp��sw��_-y�U+�\*(�xT�$O�|���xzU-W��$�A��N�aq Yf��JGXA+Ѓy�ԭCL��{6�'�N�t��Q�u�+m��|�����wH���0d-�x�&�X�?���t�˧�p ;��UQl�7��A�C�A�FX�|k@�8c ��ßr�^��l�=�u�bg0��lO�d���υ9`V��� �����+NMxw/Ei)f��'F�A$X�m�t%~̰�A&ٙ��x�d�
-��eVR���T���"e�\�
IT��⾍(������,��'R �lzr�����sx�	m��ƿ�GE=	7Ș�fT���<�3���;x�p� �晋��ܲ�/��<�O���l�a�$�I���d^K�P�T,A�}�ꤕ%c�f�o�F�-�^�qN�a�؛�vK,aj1l�檄�АH�=��[�\����q���F[�^yu��lP}W�tU�:�K�o;c������g��ib�%K��E�j�B���)�j�Q-����VU��>��r���3�l�
�ҩ��G�g�c�=U���g�^Q>q<��Sx6�L\�)B���*�E~��Ƹ�!e&r���VI[̓NAއf��t	�m��}�,nyDz%<��pi�޻�hcI��
yA��| Ύ�o�`��z~g������3�r�����`�@'�;�T��h��`#���7k�����I��&+k�4��*B#a� ~0��A3�$��_��_#����2F<�M�S��֯�'��rrm��_���M����WQ�٩����F�S�_�f��I!;ϖV3��6�An��%�1��xQ�)�P¿>��z��'�/['�SVZć�`\\�0���w��f���T�F��
�kudXo���鳍Pe�(����!�6Uw����W<�zj�����82��Nu�S���9��U�J�sy����ޮ�T� �<�&�=���Q��Q���v`'Luc�qWO�	MH�w|��	���t�hEʤ��V5�����sU�,M���K+f4<�&�꫞�gs�E���tSk��{��%
�C�Z,5*pL�BX�	VN�6Mz��A�m��G�:P�5�jn/�*�i���qO�_��h��.�φP`8�$Odj8C݊��,���^��g9��n�wʋs���Ծ�����3�ӎ4G�����i{b��4x�@��?�{��l������n�.���m��pڵ��4��]�دi�V��E��$�C!_�n &3�ש��o�$�x{i��է�_�eJ�R���}`��E֬N��}�2��Ͷ
jߗ�kd�d�����D��������+.Q�c��?�m
c�(�8v!uQ�Te���U�K��^�8p�u�>i�(˯��g��1����N{�x'��6
Mg�P�# 0�1y���w�B�1�2|�nd@Mʔj3���������l)�o����h~��z�P���Sms@���s��3��)�Uyo@����
�i�w	6#lxߞ,�'�כo���-�f�u��4y��鬕�Q�56��I�#S�e�Bc�1�O#^��m���� ��o�'.p.N/�B��৕�P�^�˱FI�&B�ē���[��Ux�y���c��G`,kz��J�*g��`����I��Jl#��$qZ�T�z|��U9�(K�6��%ΰ����b�I��P���o���<w"��HXǙ���m���k���ea��ɏU�P�W�W?��S�*�l�N��^��H��{8v�|�F�
k�S������wU4 C}(��OJi̥R��,?\�@*[�Z�V��2K������!;�tܦ��*�y�R�֭5�N����6��m9�Zw'�s�݃���Gk@Z�W�W[R���Ku�)$����%d��ȃ�2N�f�8Tۥ�/���1�*_.�ֆ���9��,d�V�:)a���Y;)�U�0��T�w�r��#2�:�Gf�*�m���S*�_����9m�_�IE���M0��f�4()��3�q�s�pu2����u�Ub@���s�R����3;���N%'MG�Sl:E���܉�p���1��9o�
��Y�Mӽ���A]6�a'T1L�V��b �I��w&�$������Ѷ� 2��������u<s��AK�$�̈́l*��r;Q1�)�&�)I�mk��K����m0�S�d�{h��D1I[n���L�o�y5j��Ռ�9o�-���&�SE��.)/�gNIwj�3�:�S~��5��z�[�0�E��-�zZIUh��Q[IE&���W��� /���l|�+B5M*C'��A�Ʈ�ZRˁI�E�N�;�Ïܐ�Z���h:K�P��L�&���O�K��S�X-Цs��hٗ���
�h �F�F����P�w���D��	�B�Kt�\Z�y$�I��O@)����V)�Ԕ��|����#�$�^�I/5-��/�R�.X8H�8���U/�pQҥ4."m��M�j森�e�kյ�,����O��M4��������7]OY�p�M��>:D�@��7(���+V%ᚂ}ڼQÙ�\!uI��ΰZJ��a��\U�cYu�>"S^�/Ւ��8�A�j���\�!���h� H���6}�o��^ԓ��vQ��@|w��>�Fw�Q�s[���g߫��}Y�<w�Q��`f��*��n�Q��F�z���4[D�� ��dapN��T����yQ
�NQ<�S?���p�C\C���&Q!�/hq�9a�Q'���GAs[x5&t�>s*��'��>�ĻTAε�|܂J�V{pK6���v\��p�97����T Ȗ��O
�� �J�I5���}4�@ID��%���!Mt�ƿK�P��b'���X�a�5(s�5y��;�}�����y�3���Kk�;+m�!�
�Z�FKM'�n{Y��"�Jd�5ˋ@�����X�϶3�N!�>h���q�!�R*�"��� �n���,�>��~7r�	�����
L1��m�����Ca�M�*��;I���TR��5��n#�R0�w�M�꾸�|
��b;�<O�}�����CJ7�Sb�zG �Ӛ�~Z,J�l�M���,���hPDB�j�����i_�f��l�!�2��eV^pF��f�U�;m\K�Y=l��@���I_�aH"�>4�-�O]�;'Z��rSW;�!�;����e8˩���N�3O�?��y��4�TnX*��⵿A��9 �s�f�x��^_�/��ъ��׻e>1
7Wũ*��M���b�@��,'L\��	]��I͋���22�h�ʞ��bNqrֶ����q��Dw���F�٢?�{�F�Rj �v��$�,Cu��ա�tܗ'5u*{q�6C����c�X ��t����+�>���R�b�j�BzR��Sco�����M�UD��B����o]2����t��S�*��b6>^,�\z�8B�4���D�]=w^���J�
j�܅#�����W��(C4�()ע hAEV-;�e������/PΥ�:a���^,*��k��H�twl�x[!��%�]|�u*�^�g�z�_Kk,x7����
{j��$�6��k��w�DC.U�@�%,Zd3���"�Ū�g 湄o��~l��@)����q���Q{�5�r��{�V�
01\f�n�vn��>|8_7N���=��#��F=|GˇF4ؼ���z��[��D�P�Ŏ����<kV�P�R3
F�GK�9h�<I��Ș�#F�W�G��Y����:�>�5�@��Z���I�U�Ŋ�#L��H|&]8�њ�z����9HձE����a
�$x�i����w�-�䇩!Z���I��x�ؒȦ4H���� \W�};������ƌ��\c8j9��a�6!�D~�]H�0�Q��y�+4���a)?��k�6zh>Wt�}+�ڦO��A���ೝ��F�X���?k�j{8�ub�vU�B��f���Be�js��EG�������m��/�Ԣ���YK�)L�Fz5�>�-��$�ے���t���4a�!M�7E�?�Iy������i4��%�N֜I�9�9y����o'�]M-ُ�q̯�����ʪ�^��z����Z�[�E5�R �&>��.�V��~�<'���o����ߗr\]�>E�o���Y�>l�K?(
\�&�5ǈ�`K��M;�ݩ]a�Y=Z�dqf2���Bc:�	�57�PN>��e-ey#l���k�����SC�i@� @�U"5��ց��<m�u��q+ȵ&laae<ڻy�6:����F^I�Û���S�h��yM����t�"�N�U� ����/6[v�xW��������%;��="��8w��SCWD{�����x׭�8��WIh��`���ie��VQ��\��I�h��J����q�Uє�(��y��J��oDPX�Q���؜H�Ѝmtd��2�Q�ڮ�A���(q?3�P����[��$d��1���b����sx@n�"W1F	rVo���w@kr�T�y���i�㌶g-_&DH�{���h�νvCe�x�}k����g�&�/LN:# �[f�m�ټ���}f"�L��=���M��a9@/���9��	ĪP��ہw�T�D���1��%���xNC�IZ;� �ī��k&⢝'�8N�������1�|�7H��b�T�ӵ�������� �̞o^(�_۬��s�]=#�]0�3u�+�K��z��+q<�O��Ѡ�:Y8^|�B����[UL���
���1�%\|�eRg&{�,``-������h�*iD���f�D��8p8����bk��)x�1Q�$��U�����j��`62L�m����XĴ[)7����A��w��~���qٟУ?�����uѣ���1n�sT!��F!�F)��i6�M��~�)�c��89�#Z��z�n�;[Y�5���5�}���Ժy��v�Չ��jm�|�kRHDjR�1�eM)q��'��4/>�#������:�N�]n�m��G%�L�\��A��K9W��p�9�p�\wU�w8BEM�❗�]���U`�4^�=����#a�OaX��'YH3�����7p�s/��?��Nrd��6���Z+�>���,r'[s``�Z�X�t3�ܝy:[�?rh3�:HP��
��;p#
�����'���J�R��(C�,��F����Z�F��M$~��W�s=Ac}��C���-q��B��+�����ȓo�ц��Oy��Y:��H�gk���p.X����0wR�A�b�����9��W�n"8�%m��qU�Z��Ԡ3�_j�Y2�!��k��r��3�u}��}U���\����d��F���6fE�	s���&����m�].��M ������HDVg=��~ܺϩظ�+ d�˪�����B@~��K��@~��ÿ��7�4��*��'&�M�gv2}�L����Dr��,�l�(���F��4Bd��F�\B�mr���Ń�=vO����n��Ee~���Fw�>�����L�,�Ű��9���'Q�_Q�ͼ��@wf�>RdY0��U�r�<ꛓ�mY�r:9�a�+^&��@\��g�]�|���r��]�%�:D���klB���d� P)ٮ��ڼ��v� ��/A��l�Ҭ�7�����ɩϙ�"�}��r8�<�V/jA�IӁ��Ka�J�R���MO�[�dx<�Al����Tn����^����IÚ�����wh�Lb�S\dB�uE.�;!�1_I�_�b��j|�f�����)� t=V`!.�'�r�~f�߮�,Ohg~����߮��Q�w�^j��`����C�y'���Am$�D�,�@����1?&�?���Ȇ�"p�V~�/��rpa��(��\��<>zb��t9��]���h:�	9�y۞�qK�tf�@�<���x���Pn�!Mpĩfg�4#�g7�q�y��7K`1/|]ݛ<�	J�j�tk��]���J�]�_!�4$��m�5Cw
�#�?����*�������z�!�~�a���H}	���E��s�Os���}�a�&���L_<�8�V�|g����P럘;
Į����Da;�k��Q�5
�i��T)�0 F��v�I�o>��<A6�P�{n^��$q��Qݲ*m|U�0j?���?�����P���;���f�� O#�f/�1>�s�Ro�.$�0@�f'�(�0%-^g���8ϭ���R���E�WKlT1^�|C���-��2�|��1��W�^dr��'z9π��Щ>|�_D��r&��d[��*��❰a�l�|�d���JKyZ�J�t�0b�$X����\S_�� )7\Gサ�5��[$.(q��KmNpH��+wܗ��#C[-�-=�����A�w�?����6;��8��.l݋tp��]=K,,v��� ���v�kD����HXV�@�o����-<H��\Dh<�*/��R͇w�J����I��n�z���D�^�Yx����(�q(�rs������_g�p��H�!��{F������~��v��n���ʰ�U�c�ݩ7����}ڒ]���A��H��_؎y|,�5Uf*ė��U����$�u]��7�t,S�=�	Ƞ� ����R�.
�����p=��@����ϲ�]!<����CKgM��~�#�p�_��Q�D
������/������B��cH��三#GO�����&�Ʌ��E���n�^��G@��KG��ڻA
��#(I�c���VM��żK�t���z�|׊����'��Z�V�ຳ�ȔO�	f5@���xݜ�#G#��7��ʮr��U��hн�����yx�ʜ�ˉv@�39E�������=7���y�G�n�O��f��X4��S�Q7ܸL�POn��N@�xU���e���
��1�e�:w�ꔱ��M@�D�����w ���޽��m�W��7���(��Q<���Δ�7�d�%}��oo�*��s)��x��u&\����t�<��kw��/�>�u����c5��&Bʯ�Fz4�U>О��`��;
M%jN�q��w�7�%�'A%gQ�w;�W�C��4MdlZ�r�0Dq�|��$�1XT=tPJ��2�Ǳ�ƺ�S���p��6���bE����ܖ�&�Y�	V�5L�ܶ.f3Ɂ�}���k��=G�ߑ��q_�o��p$�BZ�B5�iܭ�m.L=~��5�V�*�k6u�ö��p�����#����*�����*KbSW�H��t����F�;=�����T3����^�$ٰt/� g]Ƅ�����?�t3�s�'��E����nDJ`��ujHzR�c/ԧ������/�L����]�`"���GI������Pf�|]Q«Kh�!����hJ%��0t� $*�ᒙ�b!��#�C���7�^>0N�73��J�6�<xE���>H� �i��D²Gϳ�wŷ�EcN��A���̀� �������g�O�w���&��I�\m��%|13�l$y���t��L�$Ns��7�b�vh�IN��H��QNIc��հw.�j$Ձ��%ȸK���3WZ��o�m>�L�
�9 �`����%�VT����R%�ؤ����DJ��T
́��Np�Gg@3��7B�y4���C0�ɡ���=Ԡf��ު�B4�y��Ž�ܛ�!"OQM�nr��u����Ci�ߙ:>��t=9�r�(��-ϝI��80��Ѷ�<��R�>z���;C��&k]D_��d�	ԝ(�7��֕<�8��1��i��lB}��`��2Vx�PV�z�Ye��o�%���ZyP����4y���e�\�t���O�x:^um����k�Fp���E�J/�i{�W���F8Y<��C��D/֗�#<ò�Y
B�Zm�J�+`�㣻�����K�|];X�ܼ�Ɔ=?ځ]�H��_j�D<�jB��
� O'W.��l��E͛~��k�|��U*�ןێ���O~��zYZ=��E��n�vVa��F�8��;��b�&�_xR�����^��35�5�>�arq��,������+�+��6r����%�f�D��O���y�1P����~����Z�	`[�K�I�OoS&-	��ځ�E�1�a�d�w�Q��]U�1$է�VuдY�7FL_8;��_��$�y��R�l�2]��vKU�K͎��@ �i�N-��
H����Ի��~5X~�(2���t�t���O���bb@������/�{.���'��G����T(l�EE��#0����g������yB�!
�#l9�1䋊WZ
J�n;��^X��0X��)�Q [��-Z�T*-à�]Vl�5�P� ��l
�1_[�lЄF؂�����Ć�ڣb+@��C�J���`I>�H�=D�
��ҫ��"�K1aB��C���2r���X�J֣S([��Pd��v0>J{a��%杍N���d�L���وy�@w���*dA s���_2˫��mȈʫ�x28��� =���a���lX~v�爧&f<�#yVoWTĆ�����i��}�D��1i�]�֫��>D �d×���<�|�NO�;��Gi9f�Q��a��$�,ړ:�" �w��& ؚ#g��g<��pN��=l�����߃���C�rw��}��3-6�=�gc���C��4QoD·e,�S���)HL}��suښ�I��𵯡Zп�����D�H�&������F�"�)P�#�͝f��4����ɚ"�~!3����{p^���M���y��XO�%�?�M�������b9�
y�{?'�@&7� �Ϡ	���8̯S��Ff?y3H��8���D�#�Z]�3��y��Q1��S>������L�w�W�'������͜�nS�E<��y7�8,b�XNq�ݿ������� -�^ؼυq.,b��}6�,݇�P�7��9�� " ��G�T��]�eнK���\���#����W�ԝ*vǘ.��!
)�4$�1��,(�v*j�k��n-H��TȂT���7�SH�_ڦ��|�gO�B��"�\W�CF=v0�& ���6KU$��`���=3v��i�Ŋ�W�Q�������h��`7�֑���9Ju`Yv�vH�ÂE��i�	=�DK�nk2���c-b�mIg���XJ�S �|��KMb��#Lk�6�ۏ-�Q����3`�w?�T���dǠbg�}I��8���v��c\f�&����H �;=W+�e�S���N1/�+:#қ�}9`��Tk7���f�'�4eO��O9�YI�ʍ���OY-��^X��G�>�dm��z���������M�٫W��j��
�@7*�i�����q�,�ۗ>ɠt��'��y�w��t���|�4YF$�y��M	�U�=�9��EZn����tss\���һ���=0��������U���V���.��a����Hm�eq����b
$��Qp.�Uȋf��_{w;xz���?��C�P�ůd>��#�6�|ik�0�핧R��#���}I����r�v���{��{�����K�`o����!�{�����aXD�xY�����! �2(��s���G7�n�(J+����n�$_���8N�[�>��}����d�m���@��:�]C���	�!;g���
\�m���aM���;�~G�4� 'ۑ0���"��N�	q"�ಲ7���P�a /mN��'=.�7�+-C��I]�TP�e��8�PR�!,�/&�w�{�Z�
�j�N�xf��h�v��ΑSY�9�����Moɳ=S�'���L��J���1#�[��'R��M	����C�IWU?�0�uY�!��Ker��=�h|�^b�|ֺD�;u�x�F_Cj��D(�d[`&2ҵ��w����`q Ri߲�Lbd7_{��X�y��-���oWeA2e�a�:�P�%�pJ&��f*����<Ŗʾxa̳[���W��z�r��M��p��ř��&���_��ؗU�5az�*\��s=��k����7���[ ;$O<c��+j�j2�!������p�+x�iVH�h�AloJ�F��B5qE�x�R�nU�l�s�µ�'OZ���U�?�~����~h>lܸ��s���l4�HB |�t���h�n9�>�\w7�0�.&��1=��WP��E�6�ҕ���I�l�C�
%Ut����bz���!�K�@?(��[�ٺ���I�O��`����X���NX-O}6E�$�kh�����u#�YE������Q�a�*W���k���؏�h���{=�(<th��.�鋕)�6y*ݪq��/C�r��
�����z��Kf��he�7�2��^�[��ڸgbq79;ۃ�.=���C9�����6
�j���#+\��p�%e>�7�O������B�^,M��B54�
 ^�94���"�`6�h�6��Zߨ"��v����Ơ�%���td��CW_�Q�{�^]X&�'o]�Z��*3��:=AlՎ)����V�n�1���_-�T|�F�d��"�Ԥ ��N�զ��ŬE�F�wvC.yf��ۆ�uN���dn�3w͍�[���G'���\�W�F&�af�<_r��]�Vc��VX��˖��@6�,�Of���7�"��AA
�������$����q����D�D��㶓�]٘cm��킁cvr�5D�V���0پ�k���!+�(49��J��?��Nf��͸4��t�z�w��?a�s���̀��G�R����l�Kf��I����S�U,�Z��$��;�8)�7e`;�!���>�?���s�ԇ����`�ђ�nٯ�>���4�@gX��fE�5�2��uu
�D�G�tX���ĕ5��=�;x��(����^Vg�ƢШ��V'�$�!7��i�s�o�'J��s��4�'�}����E�R���-�ToW?Y�,M�� $�c����ъ1��o`�GLԅ��>�L��ρ2�̘j���ެ�����1���vRN��a��Ū�f���Y�g?S�������	S�i�)q�,ߟ�sّ�r�#�P~� ��]��/��i�ci�Z3%��|k���F;��`����"�.���-���w]<��!�=���hF�5�2I��!��oA[yX�4�G�C̙�#$]zc+�8�sO����c�G�a��P��m��,ElR�aĒL���i�ۆ���D�9���B���ᵡ.}�v"!��r��b7�%;��������( 1��m�v�1it<V��B�� �p��v%_��O�K�>������v�c<��b!�ͪ}�9��<��(�
����g9�;P�j�� �T�(}NwQO��h�L�����ȶ�F�6\s5�|�O������.�к�4�w��2����'(j�����z�g(��������L���r���f(6C�AM�GYb���Բ�4[禊��&ْg�#k���@�f���Y�eF��g��ڝ�Az��t��U;��s!{�l��밪K�U�Dz6o�*��CEkן�sʞN���e^r�<�;��e[u�ړ�EÖ��sG��?����ݔˇ[���s��-n����_��~7�=��O�kk/U�-~|���э�â>gc���p	��5���ߧE�$" g��j��;�t��79ܸ �P�6�'-�E���u����$�ҡ�8���>�oƒ����E�Კ��9��;��^��O��,��Sq�aɕx�����Ԭ.�TPN�ם�'��O*���A�5��� ��+h":P��!�s�b�,��5�@��+��Y.o�.�O�z��3T@�����>��)¼b�*�.D�ݯ~X(�8��l��,y���Rm�2�d�����vBKo�B��V��Χ��H��Z1�_9�k� +�ʟl5JA
:xXt+Q�({�@�4Ļ�)Ǵ���{�px�%tj�&۲\c�1��'s�*Z[���4���(V�Z�]xq��$�:9Wi��sKm1<�Nnd�ߧVG�j�qm������7�0�ٴ��m�AK^�v�)&�FK����A+�Va: (���5}�x�}���6�qz�${Q���C�_#t��7�]� &m4�Ұ���GT7���=�X���D�?;�A#/��;ȓ�ze{�Qˎ���.����}d�C��3�c�Dw�v�"~�_�1���H����r�]�F�n�!$��X.��'}�3����&Y��5���JZ{��6>��I�r�&����N��O#�'x*����}�} �}�ԉ���]$����Bnq�<�`+l�Dϧ� ��/Y&D��(���d��nR�a�U)����+d��1�q�̺��l��"A}i��n(�3���H3\�M�@�Em0{�)xɅj
ro�-�𻩧�q����F泸u�"Qkpy�I���.ѹ����3���&���5u6���F��a�`���\�n�"�eiM��&�b�����g�ω�G6�n�d��^^��Z����65G��A�#)Nź6���F�����k�,G_E�L��Edw��,/�}(�d����Gh��b����CN+_ y�D�Y�M>IcT��s�޻���86K�t0ӵ����0q(V��s1Vl+�m�g^��w�Õ*�slm�k��C�!Ҁԥ�爘��W,=���!�Ǔer��԰�o��[�!�_��$�,��c�=�К�^��G;��g!3���I��I�J��L�e!l�E����s�K�) w�b!&!����W��rC(_�d�Y ^�S���09
:{�9eW�o��a7���|��~�A~M�`���"�AǸZ�l8N/DEI���z��5/l�H��uW*r������[6s�b�O�zt�*��k|���K谁j�٪_�l�&����~��$���E�(
��@�����/�I<5Z�-e���� ��;ƹ_ܪt~e�b|�œE��q��΀����B��f����f�:�~���f�=�_9���	�\8�uֈ{ָ)�67*�T��G	)�E�T	��"F�5|s�\��w� �y;��=���>S-w,��W�-���
��젘�_~Pi��Iw�g4�1 �f�\��!�5.+��DO��cN��&g��sڛ����Sϻ�S�OOR����*&��Pp��`�o�T6� �o��|_#��:K����ȡ��w�� t�����G3r��AL�}�$}ԓ��
�+uYn'�Z�K�$!c�5\�(������=1���\���D�H�ğ��55�{�����}���W��=��ۂ��$u��y��b`D*�T/�'q��mAt�ŎX>�$s�D����p�hʒ41L%sm���gi64��w_��R�>0��'�bx"��� �Y�$��a��@Z� j����np�/~(b�&��4P��W��g(&w�9����Z����1�7�47i	P+��xKl��xX�b.����G��`-F����� ߱O��I��S�x YÀI�Ǝ�~���PS�Y=��_��z�<0e0��r�͒�W����ژH�,�ϱZ]%tE�ר��fF{��;S��+�����ah��M*}��F﫮S�}�x����c
�����] �5��ҵI'~�;$�,�-w�`p2p4��{ױ�`F��5�
?4Տoo����뱣g�#s��K�cb�T�3;�F����JW��ؠ�y��=.��M�$�1]�����\(�Vm���e��?o�&[N00ţ ��l?7q�#IE����l�+*�W�R���3s�D��l�8������9ϱ���X�/tV����d�4��]%�;*y:`?�����U�O���� ����� #?L}&߄��'��ݞ�08nq`F$ ����� Lg�(��S܍Xb$�U!�"1����𣯺o �j�$i\��B�m ���_��_'���?RE��S+R����ZSˌl\�/�{��P��O�Ө%�q.���89C������ZguO��(QHl��x�Z+�3�f?�ьu�ᕠ�"���a�u��}����_*4X�d��S8Uܸ�Y7���������]���i$�-J[���G��in�~��[ן"�Sg�4��\�ņR�ޢ�&�8��D0p�p�G�kh�Sh.o������A�9�a�zE����L��\=I�����S�1t7�-�8��x��L���H���z(D�陹+�u���������V~~3O��`Ym��Z@V��jjl|utI���͕�Y�Ʊv�i��T���dC��e�&�f�o��ݬ���ԑg�,�"H��ҧb�>7�3h#�}3���b�#�a����@8�#G��Yيb+��M�D�K�(�b�4�� �+�����>A����ǋ.���}����X�;a� z��v��%SPz���E�i��@U!�u��RI>O���);YB�ׄ�2�!|�ӵ�L�Ũ�%���d&��D9��<a��ca�e�@0Nr�@�qP+A�����`[���#����9�R4��S��M�hi�K/�D�A}�ݨdN8ꏑǅ��_�(c�X�-c��ȼz�рD��8cA|A���0uӣ��dW���ܣ��z')��Y�,ֹ[z��h႞�jQV����n�7�wZ��~OBL�u�a�;�������k�|��3t��4R~ ��נ*��T�^���6W�ԁI��y�}���S��dS�SQz�B��C2Mw�v���p׺�D��r\Sr�cJ�B]P�JaR�½�|���ͨ�/���t� ��4��RǍ*�n��hk��j��ģ<�\����;���n0x�qC����K�ر�%siw�W?)���-xfzz��+����a��Q������E��ӥ��b}1ӝ���6r��5!�����D�e�����L����
đ"�6f������3/�e��(���v+��\e�.�E��G�u����*�	MV�"�DN�o�
��Q1��T#�Չ]��n�G��F���#�4(�/]�v��x[�?) A���>N7�>� �țI�j)�7p4B�Ж�dUR��dӵ ���PǠ�������80����Y��~��pL(b7NO��_�'�W���A�@:��/@����燉�b���1V���� c����^%�ș=�sR)%*Tt�X>�QN���m��O$ms�WS����M����@r�����&�;%Q�@ք�	��h�i�s�5�B��C��1{[L򀣕�`�	R�����;��t�ܹ���ő��7<F� ����v�����B�9k���f<Ԁ��7�.����s-�k�g�'i�)L��B���BL,t���6��)���;�]��V�E��)��*��H(�$n��udj�����yc ဨ�xn	|��F�fۧd(բ�J$���2G����c_K9�=*ʞX1��kA[����ޣ�zf�?*�Rq�彯�o��
u�K!�T�A�_K�35��π�sW������b�6/S/?=��FJ�4H"^�*%#�gZ��	��������qӉs1�w�X��k���gB�`��[gJv&U�=�1�XV4�9��O]ksޯ5e�3�;�n�$XA&���ҭ�UR���<;��\�u6J3��5}��[z�ߓE�u*Rh8�ل8�񎻠���.��=N�`ߑ�f l�?��������:�	�X�κn�BTv5f��~�61Q���� +�XY����Va7��M�D\R6���.1wo���B^Р�ګwP�ά.v�
��́�ddN����YC� ��8#Q��H����ʏL��z�h����5�n2q�E�}�sI��{'?�kn�=�¸6��i�)����s��a��@�տ4������hѨAՊ��PL]9:5}�8�e��b_Z��0|$�>��7r=*wy�W�{G�c��,/,��"K_l��﹘��]׈�]��\��毾�J(a� `N�b�ѳt2濒��da���7�Ӽ.=
2^Ƀ�OdY�Qj_'�.��" ���)"5������ԃҦ�}�FN�����	�>+=�� FP�ѿW� ��*g���%���V��4=��6]��D��� �~<,V�N��$���5X���ٌ�2��(�F1G&=����.?a�;�m����B{�b�u��`	�q�X������D�X"C��Ա_�������YYrI�%pc��Kr�D\�goZp/���<K
%�Y�O9�$�:�F��&t�ŝ�o�\*r�#��̻�������h�U/Q�!,��b����6�e�-4�Ap͟=��� L�����i�8�)��Եh�����!�?����k	�$]r�k2��N,��W=�y1��e5�W�^����ѝ�3����G��"~n�S2�=G��T^���+����y(�G�!�ar�pt�� ~�[9��3$S�wW
z����a�����@5�I(<t~<hs��B���e�i���mߖ�Ƒl,�%7��|Y;٦�r�~�W��u)1Peoo1�o�b����0�z�K�1����U�澒|���X�X�͑�~k,V����Z���%W�6�| :�ë[�hh-C:Wj���:P�bBȇ%���6�L��^��飌���[A��b�)c�Ww�'%�� }���D*�3V�T�2�H���Cp�����(}c�~<Y]Jxj��&��G���ݜf�@��k�U�b��͞t���Aq��&�����]R%��B�x!��/3�Y�/�X�MY΂8Fѡ�o���L\o�h�([��/p*�7�-���9H���u6�^It��d4d\�B���/=խ�:B���#�� �<���G�def ��/i�+��o�h�L c�fa_�Ԉ�P����C�����4C����l�{�n������g������Ks�v<���gJЭk �>~P��y#+ע��S['ʛϞ�|3�H|QK�n�Ĺ)�Z�j�!]kġi��jUF[�rv<�i�с�����+���$V��o�!L��=jHE�Y��j����r�R�%1Gz��c׀_:�">��0E�6��\j�;*�P��"�f�+�v���6�5���p�xG��t�|H�4d��F��h�_i��i-�6�
ȎG���!��<�B U)��lHX�,R´��'�!�I���0?|�/���q��/��`���d��	��}�Zȳ�U���3�^�m�Ex&!�|�ˮ(i�+��,����3����!�ǈ��cG:�[ ���D�ڃp�7U�7U�o+�[IQ�Y���Bqd_�$��:J(-'�AY�1u��(1 ��-���I��(*&D����Os�p�ff=7�Z�[�B��^Y��&���/���Z��CG,B��?�g�_�4+���U���3dcU�_{w)Ŏ�����8A��Oe�K6T�pk�d҅3�أu>�C/���}4�i*��ׇ�	L���.4�)��	�'&"R�J&Məh�V�=��o=8BG�,FT5��W/S_[�c
Z�G��
l��J2��C���U��l@_���bU�I#ȑ��G�B�t�"'e����7��+��E��֊8[�/�̬$��*M1���:�!��M��#�����1�@�:�$os�(�W*������pf����L��u����`㸦CC~gc���ŏ3��6��O�n��& �	b�/>aFF���������%�j�s*�6��/ͷ3���g�m.�]W�Z(������Z4�H$o6�4�틣u�;a�
�[}T
����y���
��� YS�ev����v
,خ"/�j�"��C��<��X��}�J:=�8Q��d��5��X�]z�fw_p���$�~}^�&�Q���Ho�o3�At�eS+�J2r�Ds'�G]rl��F{���[fc��/���J��d�Y���Yq3�FaS���u ��Q���G3ݾ*��ř��>��@Vu
�J��K���O��qӈ/����Į�W�)�5��
��_�x8���݃�|���T�>5���������F~58y���f;�g,��A`���0�D se���%0�&'x�=���c�c���%V��A�����}�Q������<�� �K��6�(˪"�W^^�?�Y��B-KԈ�s�����
�y��Ld�f�,&?t41�tS��ʐ�R��j$CT̮v$��=����)�M�<�<픹yWW`���lR���0[K�0 �Y�F��WϾ�)���Ңr�W�dbC$�Q�Ƃ�Ҩ'r5<?���c7C�K+��U����{zcb0���р!BVW���z-b�楳�v��c�Q�ף�;���"��.�v��r�[��+�!�+t:{�������(���q�ɴ���H�UY� �����u$	ؕV��y���Ab#��Y��?��Z�b�_CuX��2��a��b�%[x�i[o?䃓�W��}��"����y�IB ��A�f<��`�Y��̦IL���-y�H[���� )Y<q�|[�(`��/.���%he��o@���p�0i�>ɮ�'�+�Lv�a���U�;Q\F-��?;j�Z��ĺF��x��k���(�"�p��o�A`��:��|C�eo�{�~֕.��qJ���2���իy<��p$�g��mE�Y��]ܬ��ݮ����/�����cL��HR��(}H�T��ϼL#�<I>,�j�K���FÛ�C{gA7\�����\�Q�R�� �\*�6S|��duUs�e�A����:zJ�yIý��#r�F�[t>��B g#i�8��u�J����*���=@���[�v�	����<3G��"��)��%=\����p�1��nխ\"�ow����䴑�`*(���Kl ��OCm1�/�+m���;�J�"������y��Kn@.���UZ��d�0��㳁Ge��G9��L`�$�q��h���/�Za�e��R��Ԙ���ra��2���E#{�Wg]�wվ����6wn�S�à�����c�I���5F��<T�i�)����(w�x�{p�:޷����f���ٶ$|���ws�v��·a
v�����o_�H�%��������-2R�(���ld�"��f|F99���9Εc�Ma��L�*��Z���o�T�ž��A}bR�rf,�b����b����r&��4��y��w"':���S�����i����o՗Qp�Ğ$��A�1T��7^�|���ݏ�a )��a� =`�rD鱭�2lV�-4��-�7@7�?Z�kg�� ��x���3���a�S˙�V8:A>%���ZR��иЦ��,��$�P�3`S8����+2ԧ���լ�}m���h)���+i��f#�����8���y���$N��RP��"�iƚ�1���\B]%�NQ$�@ϛ���.	���"|��E��$�5�Q%�[�q��X�i,�j%Mdkң��r8sfQ��Sx1�ZG�y�����"�Wvv�-��<lo9=</�e��K 3>+��+<z���4v��z	Q5���x�[�ej��4P�1x��:�y�YYd+�^�9� p-��N��}|���/�k�e.��F1:��F��ǄI�L�_��wҶK��4�,7H�K�%]'��4N���JF �8LR��+������y�Aژ��K��`(��l����#�W�<�r�CA'n##u��>���u��z�m3ppX���"f�e���-K:޹5Xu/���ܖ0��:�l#���/|k�ց��Q��I$;M�Ih�%L4Ƨl���IWo�}S�D(��GBZF8�i��c�K��� 9Om/|�WҾ�w�=DڨH�C��w��>�2�֑�I�V������'����D}��t	p[����K8Α�ӻ,�z��= -��*�ɩ����uba%`�DF���}���(����`<ں��,�D����wȗJA�n�����1#
����,8�pD��i	s@|�Z��b�K��
����c��N�S�X�9�UgP���,�^�b7�:�Q�VMbu�������"�y�n����[IB��2LPB��W�͵2��3Qp(� -��x�*�ߞ�Y_\�Lp/r��Տ�|��Q�":5X,|L�����Ԝ��tf�Qth�g���%������Glu����������F�+O�#��jeT�m�yC�������ns�1��� ���&3F����ӣU7�8s��U-7�Ǯ�^���6�������d?A�7��1��#ێ��|4:cC�{��=U���)�<�Jͅ!Lj�	��-\�!�A*�og��vNd{�;�Nd��3����3��1|�Q~�/�͕�z3���Xȑ�qT1{�$�j���j5��XФ�R��z���n�wZI�&̍\�������tr#<L���+��F�j��?�a�V<�a9����i�Z�-ne��Xh.��Ct����]d2�s6#:qk�!�XP���`�n�~��vy|��d@���k��K������2�_S6V�%����1�wEÏi��Į��O^�я���{��J�_����f���q�.k���,!/�2	�i_�Y-�+:�l���%:�o#ӝ��l�r{T�n�DU�0�����i�V�@3�j�or�y�7��ot�Prv�ҟ��v�m/��6��?�T����;�$&}yi�L,G�я��©�E��c?k�8�ȳ숤�i~Y"������v�ņ��<FN�|+,s�:��1O��k�tm���������������b9���3(hy��}����Oҩ�,��^7+�^C��P`�3Z�K���.% �����Zi���n?��	u�bо�>1�����m�R��9��*���+�`J��|� ֖�?:��C.�kp��� �<�тN)^Q�E�=k�]����^�=�C�T���*p���iIz]������&>̲��2b��i.zp�T�*c�BM��ߍ�����/[5��/�
O�i:j<4�'7���n����b��,�u�a��ERy�B	{�#s�o�MyF�l�?앨�{p���/KD��0|��
��*�����rm\�S��$EǡyQH�k�ds�:�D��:�Դ���V2��;"�/��t�h>���9����3Y��^�=/��S|�y� +Ď�M;f�$1���f@
����-����8:�������Y���(V!�j#?�B�f STo�P�|$1�t=L��qagPq�����yc�c�tu+%V6��1�q��6v \J��4�J3������������v.�!�XTꉆ{ ?vK� H�r�������̃w�]��@$
5� �t�J��FU�0P�F�vGOS�.b�޿Mu�A�T��x,W�ĳ��RKw�ʩdٳ����E�(��A�`��z�1v�%��*���~vˡ�W�,й^����Gx�1��fó�wVng
ĉ9��r��Y���� =�����^��0n���=�����0��/
�*ް<�u[aŎ��OK��v�Դ� 9�E�i�'�p�`?�8�.	�"�6���*�e��}��`z��3�oDӝ��� �5���K%�H���^��q*g�|���mw��TX6��$�<�<�6�X���l�$�Ԭ����[��n�D2�;���@�JJw��y�ўS��3���5��Wg�8�.�33�A���H��P���T�l�R��x��RJ~���(�߉���`���q��B����P4K����,���Đ_�o��* D�C0J{�q%٠L����Dbׯ��}+��t�d�U��q�W>i��&�ݘ��G�σ�F�'��Q�f`�>�s��m	�M9Uj?O.9n�a&�l:T����}C��D�$�Q����<u��]�^�]�ir��'6s���Dρz�6�?Q
�$�3K��������}�Ur�#�:�t63� ߫���h�}�أ���"y��r 1�vT�'�7�&T�æ�����;;n���a&Zj|Ԯ�	���X�V)����6:����=Ѐ�@3&1z���+煻��̈�AK:,Ƨ�< �o�|����
7��Yc�N"wn�T��G��]Όir�����fd��7Қ�QmR��lʙ]mA6L9���)�l8��:�N\�|�G��ͬ�}/F�o��rYӧ�k޿jT�v^����#�����	�����8��z�c�_��=>��Fy#Q��c������g͸�-UҘ��k�(G�1̆����1L��cX��Mƴ���Z�= ��dr$9�A�� ����!E_�[p:�Kvk狂"]s����Q�2��=��~ǭ%�S'Py4���'�F�� ����s�}���00ؘDE~�����u��>�\{%�?iZ�ѤC�=��Zs�����$�} (�r�*�C�tUXR\^��Q|����n7��j̽����O?��nI��Jۼ;B�D����s��ޑ��w�`�����9�h�ȇ∄���ޠ�X��/ �x��A��P�	t-3u_�>7�&��_�	�a�P'��B��(Ac�g�S�۸�)��O�`���I�?��ں=M�nγ7���+��_��m�҈�[��G	��y={�N
�]�Q����(���WX�CW7�O��eSsC@f�����K��.֓����U�hTOS��2^�)����2L��Aix��u`Ssv����ݱj-��jvv�8�=�,�AFV��{���^�2s6�`¡��!UmyS���Ojk���=�=�œ��l���,� D
X�Ū*!eHЍc��+ĸnS��� ych�K"�Y�u=w�}�h��?�3	i���Gɨ���!LA�˒�cg-�Y�۹���T{�V�i���pa����s(r�hm�����jðk�ڸPa:�e���� ٯ5�%����M�]�a7� � ��wgߘ�����^������i����|��;V�� �S������/��gw�U�1�gu��E�EP�6(U�sf��H
�2��~����sB�>^��J��u	��zճeSje2�~���� �
���Ů�Ef�^c[�"Gf���<M�fp�f�YqsS��ƭ����ڳ�U�m a=D, ��qJ���̫�~��iR���':/M��3)�x�/�a(?m�[ё<�8Up���M	ޱc���|�^���w���2׽E�P�ʀ~S1�	������2,[��C�"�_�0�`��P%��j�P��0Mm�M���A�m�=0�<�d)�v�� �C��O������{��N%�M�'gJ���%/���?š��ޯ�4i�w�p���(�D�����/��>n]
D�5}�a��5��W���[�$�KA�1�G�<��������>%T�m@����VR�� ����>��չU%߂��e�r���=����M��E�	���w��7E)��uQ�+��� Lȫ$d����A���t4�a6�G�������$mU\L19�7
+8�}s�Gŕ�Ӭ�ph��Zf��[`/��oU#��vi�
!��.:�����bK�s�ԏ0�P�鶡,�6_<������n������P��Ո{�q?���_�����m=��`�-��R�q`Y��9Z������%���9�����M�M�|���í֧��tO���yTߒ�m��$(�Z�A�h�\�Lj��b=��JS�Z�hB���^�����_�C��0�c�mQ��3@��z�i2MYԤ���_�Z������<�7�-�w�-&�M��h}�N��;hs����5��<wp���
?�rK!���ȗ⍵���j��� [5���B��K�K)�z]����T7�|}�� ���d��6�\���9�x��A���2�
ҬM\�7����z��75DO/V��5F�[���H mf,Us��6n]X��r�v�?����~A�W���t�)A���1Q���
+z�d}��3�Z��N�$�t��C�<j�M�O�l���8��2�6��ȟX��*e�8"$!����5	rp��1�;)ȗ�Vrբ��xG����.�����O�#�(��Eէ��՛��p�=�� ������bv��/4XX�ǉAzMu�a�t� tA�<Q��4)�8��!��գ��F��ǈ؂�Ex�R��|�׃%=��9D$-�����L �?i ��¢���H�)h�k�$s�>��HE��sc��i��;�#j`#��mP\���_V�9}�t�,54u�#�Dޜ��j/m���4O����fGA=��Ot}C?��k��'������e_�l��ON�V̜Ӄ�qC5Q�Ȥw~9Ӊ��G󛻸�a8�D\|��T�WZ'���Mғ�$
�
}>�P9XY�|�C��ݯ�J
�slm�;y��ˁ�d���Fq�bYz�'L��/N��sƚ��T5V�S�&�����?�����\��<J�������:v�y����"�4��|4,Wm1�c|�����9Ĭ�,W��C-�	2)_v�M}����;�PTEL���2B,��dΫ�"���r�D�#�aX5-h҃�CƘ�صZ�f����[|��=�k�C	�W�-2[�'pcd�&��ة�~��U��t�F��� 
T��1��I_��:842;�8^k*hɥn%~䜸Q';7q\NW�cPS]}���V}���ͣ�Zz�nz���M��Qs@�Aw?����(ǚ�e|�'�lrv�?"�"�ЮC���#i��K�-6�5�{EC��/���F3�ŠU�¶ɼ]�T��T�T��Ck�l��\�>l+OU�Q7F&�.��E5���y�� ��Cq���EsRuk��4LFPҿ�"�m���PE.�as�Uά�e��n�]�6$� *R
�N�,�����|��nn��~f���J=1��ֽs��="��C��7+���%�^*� �@�5�wB�8x�
T6-�����G��'d�f���x��J�j�1IXA^�ғ^�^���`xS�@.Ԫ�׸-��*Վ�F�5�u��g	�{���i�G5N�Ƨ��O��p ��4r"�޷Gr�@�d���߷�{�a�G3յ69&CD���7�����ە:��7�H��᫩
.��U���vt��.(Lw��:���ؖ���*�}ӧ0��W#���0���a�̈$�tlAu�*g����f�V5���|�T���j��� G��{�Rnd̖Ӹ?��zz����/�l�����D
��?F��������~�Bf�4N
awc�(X��7��r���R�s�io�
E�W�9���v@}��{��{o�oR��R�[E�7	�D����@Ե���D�j�{~��WjX���X��6ۆ�f/���S��t@�?��xÁ�e)a���_�8dR�_�Tɞ.�g���ex�@�^� ��X�,[�cY߇���%�c�W�f �*F�U/^�i˖�By��XZ	r<�'����%��z�Tw�^gM�Q��ʡe�����"+���n �#4��=�v��J�`������i)�I����+H�=˗'��������0� �
W�*��#�ϕ#�v�7��{��z���1t0C�u�e����` lT����<�gX���r�,p\g��[l��%N��e��1`5��7EV4�+��e[��ٞ~`9��2�����L�����8j��'�"������UrR98�b��%���H�`��� #c����JM�ń5M] ��{_ŠZKK������Z��ĵ�`/K��KeD��8*���:�S��K?��_��N��R%͏��O���3���^�kf�����X�g��ִ�Ӫ5�v!�k�|��Kv�+���I������5町��ٻ(4H�U�v�o��9wV[�f%�+�ó&��	�I���J�A�o��m$����p�`��t�<0Jt識�e��Ig!�|�ӥ����վ2Zܟ��tV;bC);۩�myn]><���n���V������r`�v9%?�؃^�a���~���p*e4$dR�<�-f,7�|d
eîV��z4�&�~�� >�V��C*����>��Z&]��5.�Ĭ(���?�i��!5e
�?�M�_lSk��=RiȲw�2Ԁ]�b�<��̋^�W�ѻ'*f �<�����^�Ha����,�:�>�A�6����)� p�]s"���Y0�o��02�B^��Mg0����G	&�ȕ6^�����0}��^&�ވ&N(c-��$�=��v�rхu���W�/t��VK����V���j�O��M�"��ɧr8k���̚;����0t�2W��)y�߈"uY=� �MtAz}�/���+�`�̵a~	���o�w���qsˇu�|�T�A�̤3}5t��4������D�qN�F<P��+���o�����<:��[2a���$������-���]�n�0�z�kx��y7J׺�5�V���|�v�����е���{�1?#*.��>� "HxN��J �'��Wu<v�8�S?�"�Nd�}�y�eG��i�R9�j���l��l��勒�O1H�`�@�UA�e[U��"WSz�{���`��Y,���R��?�t��*����~1����B1�ot��e]��t�
�& �3�"9��HNW��i^�]sԁ�gP�$�����f�J��J�I{��o�&If�>�;�5�4��Sv:�����U��3N�3ӕ(�4Ug)�O-�9u g:7tY��/���eLX1��ؠ/ɩw#�Z����4��`��l�T굾�T���5;̍����b	>va�� �p�vw� !�#�X��NŘ��K������}��� n�7�F�,፻u��F�1�����$!���;+x9�݊�	oWS=r?�6�E@�r�Sb����җӣE�M���t��������G���^|�Rp8Q0s��z���%"�B���}`F%�:S0T������|�^4�p'K+����ݶ�źE����E�ZT��WK�$$�����gK��\I[�G��Z���>�aK�X�`0��D�Q��nc4�P����|5:���I=���(nZQ��K�̈��ќe���
�ҩ��x5��#���,�J��n`e��[=��k«��\F��n�1-ﺅ�
WW�Et�nDj��Kh� �~2��7�@������^c�~�o�:,5zL�[���x��`?�-$�e�&��c$�����
����V��:�6���N	�P֗E�W����do��̊xw��O���Q��Q'�O����o��z�����Dr0���Hџ���p�d��<sފ?�����]ns@��l�^[\:�a_za�m+t��_j�����¸�Z|����p�S~lP0)�&��í��)�"�P���*�'�Lֵ�w�nv�ѷ��9j��8�~	����R��x�96����Q����De��U(�O��Z��F)���Uqfo+4*;����������>�7��������1O|��YҮ;es��2�[�\�������	:e���,��pl�`��9��ɦ��	���������
�J��@J]$�ڡ|*h����K�V��r3j�Q��;"1	O�K�