// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 15.0.0 Build 145 04/22/2015 SJ Web Edition"

// DATE "12/08/2015 00:10:57"

// 
// Device: Altera EP4CGX150DF31C7 Package FBGA896
// 

// 
// This greybox netlist file is for third party Synthesis Tools
// for timing and resource estimation only.
// 


module ifft_8p (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	clk,
	reset_n,
	sink_valid,
	sink_ready,
	sink_error,
	sink_sop,
	sink_eop,
	sink_real,
	sink_imag,
	fftpts_in,
	inverse,
	source_valid,
	source_ready,
	source_error,
	source_sop,
	source_eop,
	source_real,
	source_imag,
	fftpts_out)/* synthesis synthesis_greybox=1 */;
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	clk;
input 	reset_n;
input 	sink_valid;
output 	sink_ready;
input 	[1:0] sink_error;
input 	sink_sop;
input 	sink_eop;
input 	[7:0] sink_real;
input 	[7:0] sink_imag;
input 	[3:0] fftpts_in;
input 	[0:0] inverse;
output 	source_valid;
input 	source_ready;
output 	[1:0] source_error;
output 	source_sop;
output 	source_eop;
output 	[7:0] source_real;
output 	[7:0] source_imag;
output 	[3:0] fftpts_out;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|entering_s5_state~0_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|state.IDLE~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[0]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[1]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal0~0_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[2]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[1]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[0]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[3]~q ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal1~2_combout ;
wire \fft_ii_0|source_real[0]~combout ;
wire \fft_ii_0|source_real[1]~combout ;
wire \fft_ii_0|source_real[2]~combout ;
wire \fft_ii_0|source_real[3]~combout ;
wire \fft_ii_0|source_real[4]~combout ;
wire \fft_ii_0|source_real[5]~combout ;
wire \fft_ii_0|source_real[6]~combout ;
wire \fft_ii_0|source_real[7]~combout ;
wire \fft_ii_0|source_imag[0]~combout ;
wire \fft_ii_0|source_imag[1]~combout ;
wire \fft_ii_0|source_imag[2]~combout ;
wire \fft_ii_0|source_imag[3]~combout ;
wire \fft_ii_0|source_imag[4]~combout ;
wire \fft_ii_0|source_imag[5]~combout ;
wire \fft_ii_0|source_imag[6]~combout ;
wire \fft_ii_0|source_imag[7]~combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ;
wire \sink_valid~input_o ;
wire \sink_sop~input_o ;
wire \fftpts_in[0]~input_o ;
wire \fftpts_in[1]~input_o ;
wire \fftpts_in[2]~input_o ;
wire \fftpts_in[3]~input_o ;
wire \clk~input_o ;
wire \reset_n~input_o ;
wire \source_ready~input_o ;
wire \sink_error[0]~input_o ;
wire \sink_error[1]~input_o ;
wire \sink_eop~input_o ;
wire \sink_imag[0]~input_o ;
wire \sink_real[0]~input_o ;
wire \inverse[0]~input_o ;
wire \sink_imag[1]~input_o ;
wire \sink_real[1]~input_o ;
wire \sink_imag[2]~input_o ;
wire \sink_real[2]~input_o ;
wire \sink_imag[3]~input_o ;
wire \sink_real[3]~input_o ;
wire \sink_imag[4]~input_o ;
wire \sink_real[4]~input_o ;
wire \sink_imag[5]~input_o ;
wire \sink_real[5]~input_o ;
wire \sink_imag[6]~input_o ;
wire \sink_real[6]~input_o ;
wire \sink_imag[7]~input_o ;
wire \sink_real[7]~input_o ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TCKUTAP ;
wire \altera_internal_jtag~TDIUTAP ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ;
wire \~GND~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ;
wire \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ;
wire \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ;
wire \nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ;
wire \nabboc|pzdyqx_impl_inst|process_0~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ;
wire \nabboc|pzdyqx_impl_inst|NJQG9082~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~1_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ;
wire \nabboc|pzdyqx_impl_inst|AMGP4450~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ;
wire \nabboc|pzdyqx_impl_inst|Equal2~0_combout ;
wire \nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2_combout ;
wire \nabboc|pzdyqx_impl_inst|comb~0_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ;
wire \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ;
wire \nabboc|pzdyqx_impl_inst|dr_scan~combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ;
wire \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~0_combout ;
wire \nabboc|pzdyqx_impl_inst|KNOR6738~q ;
wire \nabboc|pzdyqx_impl_inst|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ;
wire \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;


ifft_8p_ifft_8p_fft_ii_0 fft_ii_0(
	.entering_s5_state(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|entering_s5_state~0_combout ),
	.stateIDLE(\fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|state.IDLE~q ),
	.out_error_s_0(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[0]~q ),
	.out_error_s_1(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[1]~q ),
	.Equal0(\fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal0~0_combout ),
	.curr_blk_s_2(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[2]~q ),
	.curr_blk_s_1(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[1]~q ),
	.curr_blk_s_0(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[0]~q ),
	.curr_blk_s_3(\fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[3]~q ),
	.Equal1(\fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal1~2_combout ),
	.source_real_0(\fft_ii_0|source_real[0]~combout ),
	.source_real_1(\fft_ii_0|source_real[1]~combout ),
	.source_real_2(\fft_ii_0|source_real[2]~combout ),
	.source_real_3(\fft_ii_0|source_real[3]~combout ),
	.source_real_4(\fft_ii_0|source_real[4]~combout ),
	.source_real_5(\fft_ii_0|source_real[5]~combout ),
	.source_real_6(\fft_ii_0|source_real[6]~combout ),
	.source_real_7(\fft_ii_0|source_real[7]~combout ),
	.source_imag_0(\fft_ii_0|source_imag[0]~combout ),
	.source_imag_1(\fft_ii_0|source_imag[1]~combout ),
	.source_imag_2(\fft_ii_0|source_imag[2]~combout ),
	.source_imag_3(\fft_ii_0|source_imag[3]~combout ),
	.source_imag_4(\fft_ii_0|source_imag[4]~combout ),
	.source_imag_5(\fft_ii_0|source_imag[5]~combout ),
	.source_imag_6(\fft_ii_0|source_imag[6]~combout ),
	.source_imag_7(\fft_ii_0|source_imag[7]~combout ),
	.GND_port(\~GND~combout ),
	.NJQG9082(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.sink_valid(\sink_valid~input_o ),
	.sink_sop(\sink_sop~input_o ),
	.fftpts_in_0(\fftpts_in[0]~input_o ),
	.fftpts_in_1(\fftpts_in[1]~input_o ),
	.fftpts_in_2(\fftpts_in[2]~input_o ),
	.fftpts_in_3(\fftpts_in[3]~input_o ),
	.clk(\clk~input_o ),
	.reset_n(\reset_n~input_o ),
	.source_ready(\source_ready~input_o ),
	.sink_error_0(\sink_error[0]~input_o ),
	.sink_error_1(\sink_error[1]~input_o ),
	.sink_eop(\sink_eop~input_o ),
	.sink_imag_0(\sink_imag[0]~input_o ),
	.sink_real_0(\sink_real[0]~input_o ),
	.inverse_0(\inverse[0]~input_o ),
	.sink_imag_1(\sink_imag[1]~input_o ),
	.sink_real_1(\sink_real[1]~input_o ),
	.sink_imag_2(\sink_imag[2]~input_o ),
	.sink_real_2(\sink_real[2]~input_o ),
	.sink_imag_3(\sink_imag[3]~input_o ),
	.sink_real_3(\sink_real[3]~input_o ),
	.sink_imag_4(\sink_imag[4]~input_o ),
	.sink_real_4(\sink_real[4]~input_o ),
	.sink_imag_5(\sink_imag[5]~input_o ),
	.sink_real_5(\sink_real[5]~input_o ),
	.sink_imag_6(\sink_imag[6]~input_o ),
	.sink_real_6(\sink_real[6]~input_o ),
	.sink_imag_7(\sink_imag[7]~input_o ),
	.sink_real_7(\sink_real[7]~input_o ));

assign \sink_valid~input_o  = sink_valid;

assign \sink_sop~input_o  = sink_sop;

assign \fftpts_in[0]~input_o  = fftpts_in[0];

assign \fftpts_in[1]~input_o  = fftpts_in[1];

assign \fftpts_in[2]~input_o  = fftpts_in[2];

assign \fftpts_in[3]~input_o  = fftpts_in[3];

assign \clk~input_o  = clk;

assign \reset_n~input_o  = reset_n;

assign \source_ready~input_o  = source_ready;

assign \sink_error[0]~input_o  = sink_error[0];

assign \sink_error[1]~input_o  = sink_error[1];

assign \sink_eop~input_o  = sink_eop;

assign \sink_imag[0]~input_o  = sink_imag[0];

assign \sink_real[0]~input_o  = sink_real[0];

assign \inverse[0]~input_o  = inverse[0];

assign \sink_imag[1]~input_o  = sink_imag[1];

assign \sink_real[1]~input_o  = sink_real[1];

assign \sink_imag[2]~input_o  = sink_imag[2];

assign \sink_real[2]~input_o  = sink_real[2];

assign \sink_imag[3]~input_o  = sink_imag[3];

assign \sink_real[3]~input_o  = sink_real[3];

assign \sink_imag[4]~input_o  = sink_imag[4];

assign \sink_real[4]~input_o  = sink_real[4];

assign \sink_imag[5]~input_o  = sink_imag[5];

assign \sink_real[5]~input_o  = sink_real[5];

assign \sink_imag[6]~input_o  = sink_imag[6];

assign \sink_real[6]~input_o  = sink_real[6];

assign \sink_imag[7]~input_o  = sink_imag[7];

assign \sink_real[7]~input_o  = sink_real[7];

assign sink_ready = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|entering_s5_state~0_combout ;

assign source_valid = \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|state.IDLE~q ;

assign source_error[0] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[0]~q ;

assign source_error[1] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|out_error_s[1]~q ;

assign source_sop = \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal0~0_combout ;

assign source_eop = \fft_ii_0|auk_dspip_r22sdf_top_inst|source_control_inst|Equal1~2_combout ;

assign source_real[0] = \fft_ii_0|source_real[0]~combout ;

assign source_real[1] = \fft_ii_0|source_real[1]~combout ;

assign source_real[2] = \fft_ii_0|source_real[2]~combout ;

assign source_real[3] = \fft_ii_0|source_real[3]~combout ;

assign source_real[4] = \fft_ii_0|source_real[4]~combout ;

assign source_real[5] = \fft_ii_0|source_real[5]~combout ;

assign source_real[6] = \fft_ii_0|source_real[6]~combout ;

assign source_real[7] = \fft_ii_0|source_real[7]~combout ;

assign source_imag[0] = \fft_ii_0|source_imag[0]~combout ;

assign source_imag[1] = \fft_ii_0|source_imag[1]~combout ;

assign source_imag[2] = \fft_ii_0|source_imag[2]~combout ;

assign source_imag[3] = \fft_ii_0|source_imag[3]~combout ;

assign source_imag[4] = \fft_ii_0|source_imag[4]~combout ;

assign source_imag[5] = \fft_ii_0|source_imag[5]~combout ;

assign source_imag[6] = \fft_ii_0|source_imag[6]~combout ;

assign source_imag[7] = \fft_ii_0|source_imag[7]~combout ;

assign fftpts_out[0] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[0]~q ;

assign fftpts_out[1] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[1]~q ;

assign fftpts_out[2] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[2]~q ;

assign fftpts_out[3] = \fft_ii_0|auk_dspip_r22sdf_top_inst|sink_ctrl_inst|curr_blk_s[3]~q ;

assign altera_reserved_tdo = \altera_internal_jtag~TDO ;

assign \altera_reserved_tms~input_o  = altera_reserved_tms;

assign \altera_reserved_tck~input_o  = altera_reserved_tck;

assign \altera_reserved_tdi~input_o  = altera_reserved_tdi;

cycloneiv_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[14]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .lut_mask = 16'hC33C;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|tms_cnt[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .lut_mask = 16'hFF7F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[9]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[7]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[6]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[2]~q ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[11]~q ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~GND~combout ),
	.cout());
defparam \~GND .lut_mask = 16'h0000;
defparam \~GND .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datad(\~GND~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[5]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[7]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|QXXQ6833_0~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:1:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:2:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:3:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:4:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:5:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:6:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:7:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:8:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:9:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:10:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:11:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:12:QXXQ6833_1~combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BWHK8171:13:QXXQ6833_1~combout ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_0~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_1~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_2~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_3~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_4~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_5~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 .lut_mask = 16'h5555;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 (
	.clk(!\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_6~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal12~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[12]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[13]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~2_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[14]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[15]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[16]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~4_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~3_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~5_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal3~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .lut_mask = 16'h0FF0;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[8]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal6~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal9~0_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[17]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|Equal0~1_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|JEQQ5299_7~q ),
	.d(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|BMIN0175[0]~q ),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 (
	.dataa(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|MBPH5020|DJQV8196[18]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 .lut_mask = 16'hAAAA;
defparam \nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~4_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal3~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal5~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .lut_mask = 16'h3CFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~4_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal8~0_combout ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .lut_mask = 16'h96FF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .lut_mask = 16'h7FFF;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~1_combout ),
	.datac(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~2_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 .lut_mask = 16'hFEFE;
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|Equal0~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_1 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|LRYQ7721|BMIN0175[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_1 .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|SQHZ7915_2 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|SQHZ7915_2 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|process_0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .lut_mask = 16'hEFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal3~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~9_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~13_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~14_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~10_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15 .lut_mask = 16'hFFAC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11 .lut_mask = 16'hACFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~11_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg_proc~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~0_combout ),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~0_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~1_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|jtag_ir_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_dr_scan_proc~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 (
	.dataa(\altera_internal_jtag~TMSUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[15]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .lut_mask = 16'hFAFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~1_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|process_0~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|process_0~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[2] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|NJQG9082~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|SQHZ7915_1~q ),
	.datad(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|NJQG9082~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|NJQG9082 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|NJQG9082~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|NJQG9082 .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 (
	.dataa(\nabboc|pzdyqx_impl_inst|NJQG9082~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~12_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|Equal2~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~1_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|AMGP4450~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|AMGP4450~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|AMGP4450 (
	.clk(\nabboc|pzdyqx_impl_inst|cycloneiii_BITP7563_gen_0:cycloneiii_BITP7563_gen_1|BITP7563_0~combout ),
	.d(\nabboc|pzdyqx_impl_inst|AMGP4450~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|SQHZ7915_2~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|AMGP4450 .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|AMGP4450~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg~8_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~15_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|reset_ena_reg~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~2_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .lut_mask = 16'hBF8F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_mode_reg[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|Equal0~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .lut_mask = 16'h7777;
defparam \nabboc|pzdyqx_impl_inst|Equal0~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal0~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|Equal2~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irf_reg[1][1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|Equal2~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|VKSG2550[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|Equal2~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|process_0~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|VKSG2550[1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 .lut_mask = 16'h55AA;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~1 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~3 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 .lut_mask = 16'h5AAF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~5 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ),
	.cout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 .lut_mask = 16'h5A5F;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .lut_mask = 16'hEEEE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~6_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~7 ),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 .lut_mask = 16'h5A5A;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~0_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(gnd),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .lut_mask = 16'hAFFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~2_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~2_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~4_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|Add0~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|Equal0~0_combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .lut_mask = 16'h6996;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028~3_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~1_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 .lut_mask = 16'hFFBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 .lut_mask = 16'h66FF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~6_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .lut_mask = 16'hEBBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~8_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~7_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1 .lut_mask = 16'hAACC;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10 (
	.dataa(gnd),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10 .lut_mask = 16'hC33C;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~9_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~10_combout ),
	.datac(gnd),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2 .lut_mask = 16'h5533;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|comb~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|comb~0 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|comb~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~2_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~1_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[3]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2] .power_up = "low";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~0_combout ),
	.asdata(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[2]~q ),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[0]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[2]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 .lut_mask = 16'hFF96;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|LCFH1028[3]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .lut_mask = 16'hBEBE;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~4_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 .lut_mask = 16'h8D8D;
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113~5_combout ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|ESUL0435|JAQF4326~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|comb~0_combout ),
	.q(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 .lut_mask = 16'hFEFF;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|dr_scan (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|splitter_nodes_receive_0[3]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|dr_scan .lut_mask = 16'hAAFF;
defparam \nabboc|pzdyqx_impl_inst|dr_scan .sum_lutc_input = "datac";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[11]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[12]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[10]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[11]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[9]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[10]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[8]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[9]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[7]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[6]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[7]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[5]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[6]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[5]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[3]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[2]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[1]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|LRYQ7721|DJQV8196[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 .lut_mask = 16'hEFFE;
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.q(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0] .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~0 (
	.dataa(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.datac(\nabboc|pzdyqx_impl_inst|ESUL0435|YROJ4113[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|TPOO7242|HENC6638[0]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .lut_mask = 16'hFFFE;
defparam \nabboc|pzdyqx_impl_inst|tdo~0 .sum_lutc_input = "datac";

dffeas \nabboc|pzdyqx_impl_inst|KNOR6738 (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(!\nabboc|pzdyqx_impl_inst|dr_scan~combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.prn(vcc));
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .is_wysiwyg = "true";
defparam \nabboc|pzdyqx_impl_inst|KNOR6738 .power_up = "low";

cycloneiv_lcell_comb \nabboc|pzdyqx_impl_inst|tdo~1 (
	.dataa(\nabboc|pzdyqx_impl_inst|tdo~0_combout ),
	.datab(\nabboc|pzdyqx_impl_inst|KNOR6738~q ),
	.datac(\nabboc|pzdyqx_impl_inst|VKSG2550[0]~q ),
	.datad(\nabboc|pzdyqx_impl_inst|VKSG2550[1]~q ),
	.cin(gnd),
	.combout(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.cout());
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .lut_mask = 16'hEFFF;
defparam \nabboc|pzdyqx_impl_inst|tdo~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.datab(\nabboc|pzdyqx_impl_inst|tdo~1_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\altera_internal_jtag~TDIUTAP ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~1_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .lut_mask = 16'hEEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[0]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~10 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~14 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 .lut_mask = 16'hFFFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~6 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~8 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~11_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~12_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~5_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .lut_mask = 16'hEBBE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~7_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8 .lut_mask = 16'hFEFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~6_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[1]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~9_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .lut_mask = 16'h8BFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[1]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~11_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[2]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~4_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .lut_mask = 16'hDFFD;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|identity_contrib_shift_reg[3]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[0]~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .lut_mask = 16'h9696;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|mixer_addr_reg_internal[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .lut_mask = 16'h6996;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric_ident_writedata[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg~15_combout ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .lut_mask = 16'h0FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena (
	.dataa(gnd),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .lut_mask = 16'hFFFC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[3]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[2]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1] .power_up = "low";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[1]~q ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_proc~0_combout ),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .lut_mask = 16'hAAFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .lut_mask = 16'hEEEE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|design_hash_reg[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_minor_ver_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .lut_mask = 16'hB8FF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~0_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~1_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~2_combout ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hFFFB;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~15 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .lut_mask = 16'h5AAF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~17 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h5A5F;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .lut_mask = 16'h5A5A;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~13_combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~23_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[2]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .lut_mask = 16'h6FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~11_combout ),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[3]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .lut_mask = 16'hFFFE;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~8_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[3]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[2]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~5_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|word_counter[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[1]~13_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0] .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg|WORD_SR[0]~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .lut_mask = 16'hBFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datac(gnd),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .lut_mask = 16'hAACC;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo_bypass_reg~q ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[1]~q ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[2]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .lut_mask = 16'hFEFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~4_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~5_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[4]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .lut_mask = 16'hEFFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~3_combout ),
	.datab(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~6_combout ),
	.datac(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|irsr_reg[0]~q ),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .lut_mask = 16'h7FFF;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7 .sum_lutc_input = "datac";

dffeas \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo (
	.clk(!\altera_internal_jtag~TCKUTAP ),
	.d(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~7_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[8]~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|hub_info_reg_ena~0_combout ),
	.q(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.prn(vcc));
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .is_wysiwyg = "true";
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo .power_up = "low";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|tdo~_wirecell .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|clr_reg~_wirecell .sum_lutc_input = "datac";

cycloneiv_lcell_comb \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell (
	.dataa(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h5555;
defparam \auto_hub|instrumentation_fabric_with_node_gen:fabric_gen_new_way:instrumentation_fabric|alt_sld_fab|sldfabric|jtag_hub_gen:real_sld_jtag_hub|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";

endmodule

module ifft_8p_ifft_8p_fft_ii_0 (
	entering_s5_state,
	stateIDLE,
	out_error_s_0,
	out_error_s_1,
	Equal0,
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Equal1,
	source_real_0,
	source_real_1,
	source_real_2,
	source_real_3,
	source_real_4,
	source_real_5,
	source_real_6,
	source_real_7,
	source_imag_0,
	source_imag_1,
	source_imag_2,
	source_imag_3,
	source_imag_4,
	source_imag_5,
	source_imag_6,
	source_imag_7,
	GND_port,
	NJQG9082,
	sink_valid,
	sink_sop,
	fftpts_in_0,
	fftpts_in_1,
	fftpts_in_2,
	fftpts_in_3,
	clk,
	reset_n,
	source_ready,
	sink_error_0,
	sink_error_1,
	sink_eop,
	sink_imag_0,
	sink_real_0,
	inverse_0,
	sink_imag_1,
	sink_real_1,
	sink_imag_2,
	sink_real_2,
	sink_imag_3,
	sink_real_3,
	sink_imag_4,
	sink_real_4,
	sink_imag_5,
	sink_real_5,
	sink_imag_6,
	sink_real_6,
	sink_imag_7,
	sink_real_7)/* synthesis synthesis_greybox=1 */;
output 	entering_s5_state;
output 	stateIDLE;
output 	out_error_s_0;
output 	out_error_s_1;
output 	Equal0;
output 	curr_blk_s_2;
output 	curr_blk_s_1;
output 	curr_blk_s_0;
output 	curr_blk_s_3;
output 	Equal1;
output 	source_real_0;
output 	source_real_1;
output 	source_real_2;
output 	source_real_3;
output 	source_real_4;
output 	source_real_5;
output 	source_real_6;
output 	source_real_7;
output 	source_imag_0;
output 	source_imag_1;
output 	source_imag_2;
output 	source_imag_3;
output 	source_imag_4;
output 	source_imag_5;
output 	source_imag_6;
output 	source_imag_7;
input 	GND_port;
input 	NJQG9082;
input 	sink_valid;
input 	sink_sop;
input 	fftpts_in_0;
input 	fftpts_in_1;
input 	fftpts_in_2;
input 	fftpts_in_3;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_eop;
input 	sink_imag_0;
input 	sink_real_0;
input 	inverse_0;
input 	sink_imag_1;
input 	sink_real_1;
input 	sink_imag_2;
input 	sink_real_2;
input 	sink_imag_3;
input 	sink_real_3;
input 	sink_imag_4;
input 	sink_real_4;
input 	sink_imag_5;
input 	sink_real_5;
input 	sink_imag_6;
input 	sink_real_6;
input 	sink_imag_7;
input 	sink_real_7;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[0]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[1]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[2]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[3]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[4]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[5]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[6]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[7]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[8]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[9]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[10]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[11]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[12]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[13]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[14]~q ;
wire \auk_dspip_r22sdf_top_inst|source_control_inst|source_data[15]~q ;


ifft_8p_auk_dspip_r22sdf_top auk_dspip_r22sdf_top_inst(
	.entering_s5_state(entering_s5_state),
	.stateIDLE(stateIDLE),
	.out_error_s_0(out_error_s_0),
	.out_error_s_1(out_error_s_1),
	.Equal0(Equal0),
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Equal1(Equal1),
	.source_data_0(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[0]~q ),
	.source_data_1(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[1]~q ),
	.source_data_2(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[2]~q ),
	.source_data_3(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[3]~q ),
	.source_data_4(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[4]~q ),
	.source_data_5(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[5]~q ),
	.source_data_6(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[6]~q ),
	.source_data_7(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[7]~q ),
	.source_data_8(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[8]~q ),
	.source_data_9(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[9]~q ),
	.source_data_10(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[10]~q ),
	.source_data_11(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[11]~q ),
	.source_data_12(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[12]~q ),
	.source_data_13(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[13]~q ),
	.source_data_14(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[14]~q ),
	.source_data_15(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[15]~q ),
	.GND_port(GND_port),
	.sink_valid(sink_valid),
	.sink_sop(sink_sop),
	.fftpts_in({fftpts_in_3,fftpts_in_2,fftpts_in_1,fftpts_in_0}),
	.clk(clk),
	.reset_n(reset_n),
	.source_ready(source_ready),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.sink_eop(sink_eop),
	.sink_imag({sink_imag_7,sink_imag_6,sink_imag_5,sink_imag_4,sink_imag_3,sink_imag_2,sink_imag_1,sink_imag_0}),
	.sink_real({sink_real_7,sink_real_6,sink_real_5,sink_real_4,sink_real_3,sink_real_2,sink_real_1,sink_real_0}),
	.inverse(inverse_0));

cycloneiv_lcell_comb \source_real[0] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_0),
	.cout());
defparam \source_real[0] .lut_mask = 16'hAAFF;
defparam \source_real[0] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[1] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_1),
	.cout());
defparam \source_real[1] .lut_mask = 16'hAAFF;
defparam \source_real[1] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[2] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_2),
	.cout());
defparam \source_real[2] .lut_mask = 16'hAAFF;
defparam \source_real[2] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[3] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[3]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_3),
	.cout());
defparam \source_real[3] .lut_mask = 16'hAAFF;
defparam \source_real[3] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[4] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[4]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_4),
	.cout());
defparam \source_real[4] .lut_mask = 16'hAAFF;
defparam \source_real[4] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[5] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[5]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_5),
	.cout());
defparam \source_real[5] .lut_mask = 16'hAAFF;
defparam \source_real[5] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[6] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[6]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_6),
	.cout());
defparam \source_real[6] .lut_mask = 16'hAAFF;
defparam \source_real[6] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_real[7] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[7]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_real_7),
	.cout());
defparam \source_real[7] .lut_mask = 16'hAAFF;
defparam \source_real[7] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[0] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_0),
	.cout());
defparam \source_imag[0] .lut_mask = 16'hAAFF;
defparam \source_imag[0] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[1] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_1),
	.cout());
defparam \source_imag[1] .lut_mask = 16'hAAFF;
defparam \source_imag[1] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[2] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_2),
	.cout());
defparam \source_imag[2] .lut_mask = 16'hAAFF;
defparam \source_imag[2] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[3] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_3),
	.cout());
defparam \source_imag[3] .lut_mask = 16'hAAFF;
defparam \source_imag[3] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[4] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_4),
	.cout());
defparam \source_imag[4] .lut_mask = 16'hAAFF;
defparam \source_imag[4] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[5] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_5),
	.cout());
defparam \source_imag[5] .lut_mask = 16'hAAFF;
defparam \source_imag[5] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[6] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_6),
	.cout());
defparam \source_imag[6] .lut_mask = 16'hAAFF;
defparam \source_imag[6] .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_imag[7] (
	.dataa(\auk_dspip_r22sdf_top_inst|source_control_inst|source_data[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(NJQG9082),
	.cin(gnd),
	.combout(source_imag_7),
	.cout());
defparam \source_imag[7] .lut_mask = 16'hAAFF;
defparam \source_imag[7] .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_top (
	entering_s5_state,
	stateIDLE,
	out_error_s_0,
	out_error_s_1,
	Equal0,
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Equal1,
	source_data_0,
	source_data_1,
	source_data_2,
	source_data_3,
	source_data_4,
	source_data_5,
	source_data_6,
	source_data_7,
	source_data_8,
	source_data_9,
	source_data_10,
	source_data_11,
	source_data_12,
	source_data_13,
	source_data_14,
	source_data_15,
	GND_port,
	sink_valid,
	sink_sop,
	fftpts_in,
	clk,
	reset_n,
	source_ready,
	sink_error_0,
	sink_error_1,
	sink_eop,
	sink_imag,
	sink_real,
	inverse)/* synthesis synthesis_greybox=1 */;
output 	entering_s5_state;
output 	stateIDLE;
output 	out_error_s_0;
output 	out_error_s_1;
output 	Equal0;
output 	curr_blk_s_2;
output 	curr_blk_s_1;
output 	curr_blk_s_0;
output 	curr_blk_s_3;
output 	Equal1;
output 	source_data_0;
output 	source_data_1;
output 	source_data_2;
output 	source_data_3;
output 	source_data_4;
output 	source_data_5;
output 	source_data_6;
output 	source_data_7;
output 	source_data_8;
output 	source_data_9;
output 	source_data_10;
output 	source_data_11;
output 	source_data_12;
output 	source_data_13;
output 	source_data_14;
output 	source_data_15;
input 	GND_port;
input 	sink_valid;
input 	sink_sop;
input 	[3:0] fftpts_in;
input 	clk;
input 	reset_n;
input 	source_ready;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_eop;
input 	[7:0] sink_imag;
input 	[7:0] sink_real;
input 	inverse;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[8] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[9] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[10] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[11] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[12] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[13] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[14] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[15] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \source_control_inst|source_stall_s~q ;
wire \source_control_inst|Add0~0_combout ;
wire \source_control_inst|Add0~1_combout ;
wire \processing_to_end~q ;
wire \generate_bit_reverse_module:bit_reverse_inst|rd_valid_dd~q ;
wire \generate_bit_reverse_module:bit_reverse_inst|out_stall_d~q ;
wire \generate_bit_reverse_module:bit_reverse_inst|rd_enable~0_combout ;
wire \sink_ctrl_inst|curr_pwr_2_s~q ;
wire \r22sdf_core_inst|out_valid~0_combout ;
wire \sink_ctrl_inst|out_valid_s~q ;
wire \r22sdf_core_inst|ena_ctrl|out_enable~0_combout ;
wire \source_control_inst|stall_p~2_combout ;
wire \generate_bit_reverse_module:bit_reverse_inst|rd_valid~q ;
wire \sent_eop~q ;
wire \r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|processing~q ;
wire \r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|processing~q ;
wire \generate_bit_reverse_module:bit_reverse_inst|processing_while_write~q ;
wire \processing_to_end~0_combout ;
wire \processing_to_end~1_combout ;
wire \r22sdf_core_inst|out_valid~1_combout ;
wire \sink_ctrl_inst|cnt[1]~q ;
wire \sink_ctrl_inst|cnt[0]~q ;
wire \sink_ctrl_inst|cnt[2]~q ;
wire \sink_ctrl_inst|Equal1~1_combout ;
wire \r22sdf_core_inst|out_real[0]~0_combout ;
wire \r22sdf_core_inst|out_real[1]~1_combout ;
wire \r22sdf_core_inst|out_real[2]~2_combout ;
wire \r22sdf_core_inst|out_real[3]~3_combout ;
wire \r22sdf_core_inst|out_real[4]~4_combout ;
wire \r22sdf_core_inst|out_real[5]~5_combout ;
wire \r22sdf_core_inst|out_real[6]~6_combout ;
wire \r22sdf_core_inst|out_real[7]~7_combout ;
wire \r22sdf_core_inst|out_imag[0]~16_combout ;
wire \r22sdf_core_inst|out_imag[1]~17_combout ;
wire \r22sdf_core_inst|out_imag[2]~18_combout ;
wire \r22sdf_core_inst|out_imag[3]~19_combout ;
wire \r22sdf_core_inst|out_imag[4]~20_combout ;
wire \r22sdf_core_inst|out_imag[5]~21_combout ;
wire \r22sdf_core_inst|out_imag[6]~22_combout ;
wire \r22sdf_core_inst|out_imag[7]~23_combout ;
wire \sent_eop~0_combout ;
wire \sink_ctrl_inst|out_data[8]~q ;
wire \sink_ctrl_inst|out_data[0]~q ;
wire \sink_ctrl_inst|curr_inverse_s~q ;
wire \sink_ctrl_inst|out_data[9]~q ;
wire \sink_ctrl_inst|out_data[1]~q ;
wire \sink_ctrl_inst|out_data[10]~q ;
wire \sink_ctrl_inst|out_data[2]~q ;
wire \sink_ctrl_inst|out_data[11]~q ;
wire \sink_ctrl_inst|out_data[3]~q ;
wire \sink_ctrl_inst|out_data[12]~q ;
wire \sink_ctrl_inst|out_data[4]~q ;
wire \sink_ctrl_inst|out_data[13]~q ;
wire \sink_ctrl_inst|out_data[5]~q ;
wire \sink_ctrl_inst|out_data[14]~q ;
wire \sink_ctrl_inst|out_data[6]~q ;
wire \sink_ctrl_inst|out_data[15]~q ;
wire \sink_ctrl_inst|out_data[7]~q ;
wire \sink_ctrl_inst|curr_input_sel_s[0]~q ;
wire \source_control_inst|Add0~2_combout ;
wire \generate_bit_reverse_module:bit_reverse_inst|out_valid~4_combout ;
wire \generate_bit_reverse_module:bit_reverse_inst|out_valid~5_combout ;


ifft_8p_auk_dspip_bit_reverse_core \generate_bit_reverse_module:bit_reverse_inst (
	.q_b_8(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[8] ),
	.q_b_9(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[9] ),
	.q_b_10(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[10] ),
	.q_b_11(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[11] ),
	.q_b_12(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[12] ),
	.q_b_13(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[13] ),
	.q_b_14(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[14] ),
	.q_b_15(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[15] ),
	.q_b_0(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_b_1(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_b_2(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_b_3(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_b_4(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_b_5(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_b_6(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_b_7(\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.out_stall(\source_control_inst|source_stall_s~q ),
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Add0(\source_control_inst|Add0~0_combout ),
	.Add01(\source_control_inst|Add0~1_combout ),
	.rd_valid_dd1(\generate_bit_reverse_module:bit_reverse_inst|rd_valid_dd~q ),
	.out_stall_d1(\generate_bit_reverse_module:bit_reverse_inst|out_stall_d~q ),
	.rd_enable(\generate_bit_reverse_module:bit_reverse_inst|rd_enable~0_combout ),
	.out_valid(\r22sdf_core_inst|out_valid~0_combout ),
	.out_enable(\r22sdf_core_inst|ena_ctrl|out_enable~0_combout ),
	.rd_valid1(\generate_bit_reverse_module:bit_reverse_inst|rd_valid~q ),
	.processing_while_write1(\generate_bit_reverse_module:bit_reverse_inst|processing_while_write~q ),
	.out_valid1(\r22sdf_core_inst|out_valid~1_combout ),
	.out_real_0(\r22sdf_core_inst|out_real[0]~0_combout ),
	.out_real_1(\r22sdf_core_inst|out_real[1]~1_combout ),
	.out_real_2(\r22sdf_core_inst|out_real[2]~2_combout ),
	.out_real_3(\r22sdf_core_inst|out_real[3]~3_combout ),
	.out_real_4(\r22sdf_core_inst|out_real[4]~4_combout ),
	.out_real_5(\r22sdf_core_inst|out_real[5]~5_combout ),
	.out_real_6(\r22sdf_core_inst|out_real[6]~6_combout ),
	.out_real_7(\r22sdf_core_inst|out_real[7]~7_combout ),
	.out_imag_0(\r22sdf_core_inst|out_imag[0]~16_combout ),
	.out_imag_1(\r22sdf_core_inst|out_imag[1]~17_combout ),
	.out_imag_2(\r22sdf_core_inst|out_imag[2]~18_combout ),
	.out_imag_3(\r22sdf_core_inst|out_imag[3]~19_combout ),
	.out_imag_4(\r22sdf_core_inst|out_imag[4]~20_combout ),
	.out_imag_5(\r22sdf_core_inst|out_imag[5]~21_combout ),
	.out_imag_6(\r22sdf_core_inst|out_imag[6]~22_combout ),
	.out_imag_7(\r22sdf_core_inst|out_imag[7]~23_combout ),
	.out_valid2(\generate_bit_reverse_module:bit_reverse_inst|out_valid~4_combout ),
	.out_valid3(\generate_bit_reverse_module:bit_reverse_inst|out_valid~5_combout ),
	.clk(clk),
	.reset(reset_n));

ifft_8p_auk_dspip_r22sdf_core r22sdf_core_inst(
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.Add0(\source_control_inst|Add0~0_combout ),
	.Add01(\source_control_inst|Add0~1_combout ),
	.out_stall_d(\generate_bit_reverse_module:bit_reverse_inst|out_stall_d~q ),
	.curr_pwr_2_s(\sink_ctrl_inst|curr_pwr_2_s~q ),
	.out_valid(\r22sdf_core_inst|out_valid~0_combout ),
	.enable(\sink_ctrl_inst|out_valid_s~q ),
	.out_enable(\r22sdf_core_inst|ena_ctrl|out_enable~0_combout ),
	.processing(\r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|processing~q ),
	.processing1(\r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|processing~q ),
	.out_valid1(\r22sdf_core_inst|out_valid~1_combout ),
	.cnt_1(\sink_ctrl_inst|cnt[1]~q ),
	.cnt_0(\sink_ctrl_inst|cnt[0]~q ),
	.cnt_2(\sink_ctrl_inst|cnt[2]~q ),
	.in_eop(\sink_ctrl_inst|Equal1~1_combout ),
	.out_real_0(\r22sdf_core_inst|out_real[0]~0_combout ),
	.out_real_1(\r22sdf_core_inst|out_real[1]~1_combout ),
	.out_real_2(\r22sdf_core_inst|out_real[2]~2_combout ),
	.out_real_3(\r22sdf_core_inst|out_real[3]~3_combout ),
	.out_real_4(\r22sdf_core_inst|out_real[4]~4_combout ),
	.out_real_5(\r22sdf_core_inst|out_real[5]~5_combout ),
	.out_real_6(\r22sdf_core_inst|out_real[6]~6_combout ),
	.out_real_7(\r22sdf_core_inst|out_real[7]~7_combout ),
	.out_imag_0(\r22sdf_core_inst|out_imag[0]~16_combout ),
	.out_imag_1(\r22sdf_core_inst|out_imag[1]~17_combout ),
	.out_imag_2(\r22sdf_core_inst|out_imag[2]~18_combout ),
	.out_imag_3(\r22sdf_core_inst|out_imag[3]~19_combout ),
	.out_imag_4(\r22sdf_core_inst|out_imag[4]~20_combout ),
	.out_imag_5(\r22sdf_core_inst|out_imag[5]~21_combout ),
	.out_imag_6(\r22sdf_core_inst|out_imag[6]~22_combout ),
	.out_imag_7(\r22sdf_core_inst|out_imag[7]~23_combout ),
	.out_data_8(\sink_ctrl_inst|out_data[8]~q ),
	.out_data_0(\sink_ctrl_inst|out_data[0]~q ),
	.curr_inverse_s(\sink_ctrl_inst|curr_inverse_s~q ),
	.out_data_9(\sink_ctrl_inst|out_data[9]~q ),
	.out_data_1(\sink_ctrl_inst|out_data[1]~q ),
	.out_data_10(\sink_ctrl_inst|out_data[10]~q ),
	.out_data_2(\sink_ctrl_inst|out_data[2]~q ),
	.out_data_11(\sink_ctrl_inst|out_data[11]~q ),
	.out_data_3(\sink_ctrl_inst|out_data[3]~q ),
	.out_data_12(\sink_ctrl_inst|out_data[12]~q ),
	.out_data_4(\sink_ctrl_inst|out_data[4]~q ),
	.out_data_13(\sink_ctrl_inst|out_data[13]~q ),
	.out_data_5(\sink_ctrl_inst|out_data[5]~q ),
	.out_data_14(\sink_ctrl_inst|out_data[14]~q ),
	.out_data_6(\sink_ctrl_inst|out_data[6]~q ),
	.out_data_15(\sink_ctrl_inst|out_data[15]~q ),
	.out_data_7(\sink_ctrl_inst|out_data[7]~q ),
	.curr_input_sel_s_0(\sink_ctrl_inst|curr_input_sel_s[0]~q ),
	.Add02(\source_control_inst|Add0~2_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset_n));

ifft_8p_auk_dspip_avalon_streaming_block_sink sink_ctrl_inst(
	.source_stall_s(\source_control_inst|source_stall_s~q ),
	.entering_s5_state(entering_s5_state),
	.out_error_s_0(out_error_s_0),
	.out_error_s_1(out_error_s_1),
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Add0(\source_control_inst|Add0~0_combout ),
	.Add01(\source_control_inst|Add0~1_combout ),
	.processing_to_end(\processing_to_end~q ),
	.curr_pwr_2_s1(\sink_ctrl_inst|curr_pwr_2_s~q ),
	.out_valid_s1(\sink_ctrl_inst|out_valid_s~q ),
	.cnt_1(\sink_ctrl_inst|cnt[1]~q ),
	.cnt_0(\sink_ctrl_inst|cnt[0]~q ),
	.cnt_2(\sink_ctrl_inst|cnt[2]~q ),
	.Equal1(\sink_ctrl_inst|Equal1~1_combout ),
	.out_data_8(\sink_ctrl_inst|out_data[8]~q ),
	.out_data_0(\sink_ctrl_inst|out_data[0]~q ),
	.curr_inverse_s1(\sink_ctrl_inst|curr_inverse_s~q ),
	.out_data_9(\sink_ctrl_inst|out_data[9]~q ),
	.out_data_1(\sink_ctrl_inst|out_data[1]~q ),
	.out_data_10(\sink_ctrl_inst|out_data[10]~q ),
	.out_data_2(\sink_ctrl_inst|out_data[2]~q ),
	.out_data_11(\sink_ctrl_inst|out_data[11]~q ),
	.out_data_3(\sink_ctrl_inst|out_data[3]~q ),
	.out_data_12(\sink_ctrl_inst|out_data[12]~q ),
	.out_data_4(\sink_ctrl_inst|out_data[4]~q ),
	.out_data_13(\sink_ctrl_inst|out_data[13]~q ),
	.out_data_5(\sink_ctrl_inst|out_data[5]~q ),
	.out_data_14(\sink_ctrl_inst|out_data[14]~q ),
	.out_data_6(\sink_ctrl_inst|out_data[6]~q ),
	.out_data_15(\sink_ctrl_inst|out_data[15]~q ),
	.out_data_7(\sink_ctrl_inst|out_data[7]~q ),
	.curr_input_sel_s_0(\sink_ctrl_inst|curr_input_sel_s[0]~q ),
	.sink_valid(sink_valid),
	.sink_sop(sink_sop),
	.in_blk({fftpts_in[3],fftpts_in[2],fftpts_in[1],fftpts_in[0]}),
	.clk(clk),
	.reset(reset_n),
	.sink_error_0(sink_error_0),
	.sink_error_1(sink_error_1),
	.sink_eop(sink_eop),
	.in_data({sink_imag[7],sink_imag[6],sink_imag[5],sink_imag[4],sink_imag[3],sink_imag[2],sink_imag[1],sink_imag[0],sink_real[7],sink_real[6],sink_real[5],sink_real[4],sink_real[3],sink_real[2],sink_real[1],sink_real[0]}),
	.in_inverse(inverse));

ifft_8p_auk_dspip_avalon_streaming_block_source source_control_inst(
	.in_data({\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[7] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[6] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[5] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[4] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[3] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[2] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[1] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[0] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[15] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[14] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[13] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[12] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[11] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[10] ,
\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[9] ,\generate_bit_reverse_module:bit_reverse_inst|real_buf|old_ram_gen:old_ram_component|auto_generated|q_b[8] }),
	.source_stall_s1(\source_control_inst|source_stall_s~q ),
	.stateIDLE(stateIDLE),
	.Equal0(Equal0),
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Add0(\source_control_inst|Add0~0_combout ),
	.Add01(\source_control_inst|Add0~1_combout ),
	.Equal1(Equal1),
	.source_data_0(source_data_0),
	.source_data_1(source_data_1),
	.source_data_2(source_data_2),
	.source_data_3(source_data_3),
	.source_data_4(source_data_4),
	.source_data_5(source_data_5),
	.source_data_6(source_data_6),
	.source_data_7(source_data_7),
	.source_data_8(source_data_8),
	.source_data_9(source_data_9),
	.source_data_10(source_data_10),
	.source_data_11(source_data_11),
	.source_data_12(source_data_12),
	.source_data_13(source_data_13),
	.source_data_14(source_data_14),
	.source_data_15(source_data_15),
	.rd_valid_dd(\generate_bit_reverse_module:bit_reverse_inst|rd_valid_dd~q ),
	.rd_enable(\generate_bit_reverse_module:bit_reverse_inst|rd_enable~0_combout ),
	.out_valid(\r22sdf_core_inst|out_valid~0_combout ),
	.out_enable(\r22sdf_core_inst|ena_ctrl|out_enable~0_combout ),
	.stall_p(\source_control_inst|stall_p~2_combout ),
	.Add02(\source_control_inst|Add0~2_combout ),
	.out_valid1(\generate_bit_reverse_module:bit_reverse_inst|out_valid~4_combout ),
	.out_valid2(\generate_bit_reverse_module:bit_reverse_inst|out_valid~5_combout ),
	.clk(clk),
	.reset(reset_n),
	.source_ready(source_ready));

dffeas processing_to_end(
	.clk(clk),
	.d(\processing_to_end~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\processing_to_end~q ),
	.prn(vcc));
defparam processing_to_end.is_wysiwyg = "true";
defparam processing_to_end.power_up = "low";

dffeas sent_eop(
	.clk(clk),
	.d(\sent_eop~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\sent_eop~q ),
	.prn(vcc));
defparam sent_eop.is_wysiwyg = "true";
defparam sent_eop.power_up = "low";

cycloneiv_lcell_comb \processing_to_end~0 (
	.dataa(\sent_eop~q ),
	.datab(\r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|processing~q ),
	.datac(\r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|processing~q ),
	.datad(\generate_bit_reverse_module:bit_reverse_inst|processing_while_write~q ),
	.cin(gnd),
	.combout(\processing_to_end~0_combout ),
	.cout());
defparam \processing_to_end~0 .lut_mask = 16'hFFFE;
defparam \processing_to_end~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_to_end~1 (
	.dataa(\generate_bit_reverse_module:bit_reverse_inst|rd_valid~q ),
	.datab(\processing_to_end~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\processing_to_end~1_combout ),
	.cout());
defparam \processing_to_end~1 .lut_mask = 16'hEEEE;
defparam \processing_to_end~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \sent_eop~0 (
	.dataa(\sent_eop~q ),
	.datab(Equal0),
	.datac(\source_control_inst|stall_p~2_combout ),
	.datad(Equal1),
	.cin(gnd),
	.combout(\sent_eop~0_combout ),
	.cout());
defparam \sent_eop~0 .lut_mask = 16'hACFF;
defparam \sent_eop~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_avalon_streaming_block_sink (
	source_stall_s,
	entering_s5_state,
	out_error_s_0,
	out_error_s_1,
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Add0,
	Add01,
	processing_to_end,
	curr_pwr_2_s1,
	out_valid_s1,
	cnt_1,
	cnt_0,
	cnt_2,
	Equal1,
	out_data_8,
	out_data_0,
	curr_inverse_s1,
	out_data_9,
	out_data_1,
	out_data_10,
	out_data_2,
	out_data_11,
	out_data_3,
	out_data_12,
	out_data_4,
	out_data_13,
	out_data_5,
	out_data_14,
	out_data_6,
	out_data_15,
	out_data_7,
	curr_input_sel_s_0,
	sink_valid,
	sink_sop,
	in_blk,
	clk,
	reset,
	sink_error_0,
	sink_error_1,
	sink_eop,
	in_data,
	in_inverse)/* synthesis synthesis_greybox=1 */;
input 	source_stall_s;
output 	entering_s5_state;
output 	out_error_s_0;
output 	out_error_s_1;
output 	curr_blk_s_2;
output 	curr_blk_s_1;
output 	curr_blk_s_0;
output 	curr_blk_s_3;
input 	Add0;
input 	Add01;
input 	processing_to_end;
output 	curr_pwr_2_s1;
output 	out_valid_s1;
output 	cnt_1;
output 	cnt_0;
output 	cnt_2;
output 	Equal1;
output 	out_data_8;
output 	out_data_0;
output 	curr_inverse_s1;
output 	out_data_9;
output 	out_data_1;
output 	out_data_10;
output 	out_data_2;
output 	out_data_11;
output 	out_data_3;
output 	out_data_12;
output 	out_data_4;
output 	out_data_13;
output 	out_data_5;
output 	out_data_14;
output 	out_data_6;
output 	out_data_15;
output 	out_data_7;
output 	curr_input_sel_s_0;
input 	sink_valid;
input 	sink_sop;
input 	[3:0] in_blk;
input 	clk;
input 	reset;
input 	sink_error_0;
input 	sink_error_1;
input 	sink_eop;
input 	[15:0] in_data;
input 	in_inverse;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \start~q ;
wire \shunt_control~0_combout ;
wire \Equal5~0_combout ;
wire \Equal5~1_combout ;
wire \shunt_control~1_combout ;
wire \next_state~0_combout ;
wire \state~q ;
wire \in_cnt~1_combout ;
wire \out_data_p~0_combout ;
wire \in_cnt[1]~q ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \in_cnt~2_combout ;
wire \in_cnt[0]~q ;
wire \in_cnt~0_combout ;
wire \in_cnt[2]~q ;
wire \missing_sop_p~0_combout ;
wire \missing_sop_p~1_combout ;
wire \missing_sop~q ;
wire \unexpected_eop_p~0_combout ;
wire \unexpected_eop~q ;
wire \missing_eop_p~0_combout ;
wire \missing_eop~q ;
wire \out_error_s~0_combout ;
wire \out_error_s~1_combout ;
wire \blk_shunt[2]~q ;
wire \curr_blk_p~0_combout ;
wire \curr_blk_s~2_combout ;
wire \curr_blk_s[2]~7_combout ;
wire \curr_blk_s[2]~3_combout ;
wire \blk_shunt[1]~q ;
wire \curr_blk_s~4_combout ;
wire \blk_shunt[0]~q ;
wire \curr_blk_s~5_combout ;
wire \blk_shunt[3]~q ;
wire \curr_blk_s~6_combout ;
wire \in_pwr_2~combout ;
wire \pwr_2_shunt~q ;
wire \curr_pwr_2_s~0_combout ;
wire \leaving_s5_state~0_combout ;
wire \out_valid_s~0_combout ;
wire \got_sop~0_combout ;
wire \got_sop~q ;
wire \out_valid_s~1_combout ;
wire \cnt~0_combout ;
wire \cnt~1_combout ;
wire \cnt~2_combout ;
wire \Equal1~0_combout ;
wire \entering_s5_state~1_combout ;
wire \in_data_shunt[8]~q ;
wire \out_data~0_combout ;
wire \in_data_shunt[0]~q ;
wire \out_data~1_combout ;
wire \inverse_shunt~q ;
wire \curr_inverse_s~0_combout ;
wire \in_data_shunt[9]~q ;
wire \out_data~2_combout ;
wire \in_data_shunt[1]~q ;
wire \out_data~3_combout ;
wire \in_data_shunt[10]~q ;
wire \out_data~4_combout ;
wire \in_data_shunt[2]~q ;
wire \out_data~5_combout ;
wire \in_data_shunt[11]~q ;
wire \out_data~6_combout ;
wire \in_data_shunt[3]~q ;
wire \out_data~7_combout ;
wire \in_data_shunt[12]~q ;
wire \out_data~8_combout ;
wire \in_data_shunt[4]~q ;
wire \out_data~9_combout ;
wire \in_data_shunt[13]~q ;
wire \out_data~10_combout ;
wire \in_data_shunt[5]~q ;
wire \out_data~11_combout ;
wire \in_data_shunt[14]~q ;
wire \out_data~12_combout ;
wire \in_data_shunt[6]~q ;
wire \out_data~13_combout ;
wire \in_data_shunt[15]~q ;
wire \out_data~14_combout ;
wire \in_data_shunt[7]~q ;
wire \out_data~15_combout ;
wire \stg_input_sel[0]~0_combout ;
wire \input_sel_shunt[0]~q ;
wire \curr_input_sel_s~0_combout ;


cycloneiv_lcell_comb \entering_s5_state~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\state~q ),
	.datad(source_stall_s),
	.cin(gnd),
	.combout(entering_s5_state),
	.cout());
defparam \entering_s5_state~0 .lut_mask = 16'h0FFF;
defparam \entering_s5_state~0 .sum_lutc_input = "datac";

dffeas \out_error_s[0] (
	.clk(clk),
	.d(\out_error_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_error_s_0),
	.prn(vcc));
defparam \out_error_s[0] .is_wysiwyg = "true";
defparam \out_error_s[0] .power_up = "low";

dffeas \out_error_s[1] (
	.clk(clk),
	.d(\out_error_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_error_s_1),
	.prn(vcc));
defparam \out_error_s[1] .is_wysiwyg = "true";
defparam \out_error_s[1] .power_up = "low";

dffeas \curr_blk_s[2] (
	.clk(clk),
	.d(\curr_blk_s~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_blk_s_2),
	.prn(vcc));
defparam \curr_blk_s[2] .is_wysiwyg = "true";
defparam \curr_blk_s[2] .power_up = "low";

dffeas \curr_blk_s[1] (
	.clk(clk),
	.d(\curr_blk_s~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_blk_s_1),
	.prn(vcc));
defparam \curr_blk_s[1] .is_wysiwyg = "true";
defparam \curr_blk_s[1] .power_up = "low";

dffeas \curr_blk_s[0] (
	.clk(clk),
	.d(\curr_blk_s~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_blk_s_0),
	.prn(vcc));
defparam \curr_blk_s[0] .is_wysiwyg = "true";
defparam \curr_blk_s[0] .power_up = "low";

dffeas \curr_blk_s[3] (
	.clk(clk),
	.d(\curr_blk_s~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_blk_s_3),
	.prn(vcc));
defparam \curr_blk_s[3] .is_wysiwyg = "true";
defparam \curr_blk_s[3] .power_up = "low";

dffeas curr_pwr_2_s(
	.clk(clk),
	.d(\curr_pwr_2_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_pwr_2_s1),
	.prn(vcc));
defparam curr_pwr_2_s.is_wysiwyg = "true";
defparam curr_pwr_2_s.power_up = "low";

dffeas out_valid_s(
	.clk(clk),
	.d(\out_valid_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_valid_s1),
	.prn(vcc));
defparam out_valid_s.is_wysiwyg = "true";
defparam out_valid_s.power_up = "low";

dffeas \cnt[1] (
	.clk(clk),
	.d(\cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid_s1),
	.q(cnt_1),
	.prn(vcc));
defparam \cnt[1] .is_wysiwyg = "true";
defparam \cnt[1] .power_up = "low";

dffeas \cnt[0] (
	.clk(clk),
	.d(\cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid_s1),
	.q(cnt_0),
	.prn(vcc));
defparam \cnt[0] .is_wysiwyg = "true";
defparam \cnt[0] .power_up = "low";

dffeas \cnt[2] (
	.clk(clk),
	.d(\cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid_s1),
	.q(cnt_2),
	.prn(vcc));
defparam \cnt[2] .is_wysiwyg = "true";
defparam \cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Equal1~1 (
	.dataa(Add0),
	.datab(\Equal1~0_combout ),
	.datac(Add01),
	.datad(cnt_2),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hBFFB;
defparam \Equal1~1 .sum_lutc_input = "datac";

dffeas \out_data[8] (
	.clk(clk),
	.d(\out_data~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_8),
	.prn(vcc));
defparam \out_data[8] .is_wysiwyg = "true";
defparam \out_data[8] .power_up = "low";

dffeas \out_data[0] (
	.clk(clk),
	.d(\out_data~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_0),
	.prn(vcc));
defparam \out_data[0] .is_wysiwyg = "true";
defparam \out_data[0] .power_up = "low";

dffeas curr_inverse_s(
	.clk(clk),
	.d(\curr_inverse_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_inverse_s1),
	.prn(vcc));
defparam curr_inverse_s.is_wysiwyg = "true";
defparam curr_inverse_s.power_up = "low";

dffeas \out_data[9] (
	.clk(clk),
	.d(\out_data~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_9),
	.prn(vcc));
defparam \out_data[9] .is_wysiwyg = "true";
defparam \out_data[9] .power_up = "low";

dffeas \out_data[1] (
	.clk(clk),
	.d(\out_data~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_1),
	.prn(vcc));
defparam \out_data[1] .is_wysiwyg = "true";
defparam \out_data[1] .power_up = "low";

dffeas \out_data[10] (
	.clk(clk),
	.d(\out_data~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_10),
	.prn(vcc));
defparam \out_data[10] .is_wysiwyg = "true";
defparam \out_data[10] .power_up = "low";

dffeas \out_data[2] (
	.clk(clk),
	.d(\out_data~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_2),
	.prn(vcc));
defparam \out_data[2] .is_wysiwyg = "true";
defparam \out_data[2] .power_up = "low";

dffeas \out_data[11] (
	.clk(clk),
	.d(\out_data~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_11),
	.prn(vcc));
defparam \out_data[11] .is_wysiwyg = "true";
defparam \out_data[11] .power_up = "low";

dffeas \out_data[3] (
	.clk(clk),
	.d(\out_data~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_3),
	.prn(vcc));
defparam \out_data[3] .is_wysiwyg = "true";
defparam \out_data[3] .power_up = "low";

dffeas \out_data[12] (
	.clk(clk),
	.d(\out_data~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_12),
	.prn(vcc));
defparam \out_data[12] .is_wysiwyg = "true";
defparam \out_data[12] .power_up = "low";

dffeas \out_data[4] (
	.clk(clk),
	.d(\out_data~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_4),
	.prn(vcc));
defparam \out_data[4] .is_wysiwyg = "true";
defparam \out_data[4] .power_up = "low";

dffeas \out_data[13] (
	.clk(clk),
	.d(\out_data~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_13),
	.prn(vcc));
defparam \out_data[13] .is_wysiwyg = "true";
defparam \out_data[13] .power_up = "low";

dffeas \out_data[5] (
	.clk(clk),
	.d(\out_data~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_5),
	.prn(vcc));
defparam \out_data[5] .is_wysiwyg = "true";
defparam \out_data[5] .power_up = "low";

dffeas \out_data[14] (
	.clk(clk),
	.d(\out_data~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_14),
	.prn(vcc));
defparam \out_data[14] .is_wysiwyg = "true";
defparam \out_data[14] .power_up = "low";

dffeas \out_data[6] (
	.clk(clk),
	.d(\out_data~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_6),
	.prn(vcc));
defparam \out_data[6] .is_wysiwyg = "true";
defparam \out_data[6] .power_up = "low";

dffeas \out_data[15] (
	.clk(clk),
	.d(\out_data~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_15),
	.prn(vcc));
defparam \out_data[15] .is_wysiwyg = "true";
defparam \out_data[15] .power_up = "low";

dffeas \out_data[7] (
	.clk(clk),
	.d(\out_data~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_valid_s~0_combout ),
	.q(out_data_7),
	.prn(vcc));
defparam \out_data[7] .is_wysiwyg = "true";
defparam \out_data[7] .power_up = "low";

dffeas \curr_input_sel_s[0] (
	.clk(clk),
	.d(\curr_input_sel_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\curr_blk_s[2]~3_combout ),
	.q(curr_input_sel_s_0),
	.prn(vcc));
defparam \curr_input_sel_s[0] .is_wysiwyg = "true";
defparam \curr_input_sel_s[0] .power_up = "low";

dffeas start(
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid_s1),
	.q(\start~q ),
	.prn(vcc));
defparam start.is_wysiwyg = "true";
defparam start.power_up = "low";

cycloneiv_lcell_comb \shunt_control~0 (
	.dataa(processing_to_end),
	.datab(sink_valid),
	.datac(sink_sop),
	.datad(\start~q ),
	.cin(gnd),
	.combout(\shunt_control~0_combout ),
	.cout());
defparam \shunt_control~0 .lut_mask = 16'hFFFE;
defparam \shunt_control~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal5~0 (
	.dataa(curr_blk_s_1),
	.datab(curr_blk_s_0),
	.datac(in_blk[0]),
	.datad(in_blk[1]),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
defparam \Equal5~0 .lut_mask = 16'h6996;
defparam \Equal5~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal5~1 (
	.dataa(curr_blk_s_3),
	.datab(curr_blk_s_2),
	.datac(in_blk[2]),
	.datad(in_blk[3]),
	.cin(gnd),
	.combout(\Equal5~1_combout ),
	.cout());
defparam \Equal5~1 .lut_mask = 16'h6996;
defparam \Equal5~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shunt_control~1 (
	.dataa(\shunt_control~0_combout ),
	.datab(gnd),
	.datac(\Equal5~0_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\shunt_control~1_combout ),
	.cout());
defparam \shunt_control~1 .lut_mask = 16'hAFFF;
defparam \shunt_control~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \next_state~0 (
	.dataa(\state~q ),
	.datab(\shunt_control~1_combout ),
	.datac(processing_to_end),
	.datad(source_stall_s),
	.cin(gnd),
	.combout(\next_state~0_combout ),
	.cout());
defparam \next_state~0 .lut_mask = 16'hFAFC;
defparam \next_state~0 .sum_lutc_input = "datac";

dffeas state(
	.clk(clk),
	.d(\next_state~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state~q ),
	.prn(vcc));
defparam state.is_wysiwyg = "true";
defparam state.power_up = "low";

cycloneiv_lcell_comb \in_cnt~1 (
	.dataa(gnd),
	.datab(\in_cnt[0]~q ),
	.datac(\in_cnt[1]~q ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~1_combout ),
	.cout());
defparam \in_cnt~1 .lut_mask = 16'h3CFF;
defparam \in_cnt~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_data_p~0 (
	.dataa(sink_valid),
	.datab(gnd),
	.datac(\state~q ),
	.datad(source_stall_s),
	.cin(gnd),
	.combout(\out_data_p~0_combout ),
	.cout());
defparam \out_data_p~0 .lut_mask = 16'hAFFF;
defparam \out_data_p~0 .sum_lutc_input = "datac";

dffeas \in_cnt[1] (
	.clk(clk),
	.d(\in_cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data_p~0_combout ),
	.q(\in_cnt[1]~q ),
	.prn(vcc));
defparam \in_cnt[1] .is_wysiwyg = "true";
defparam \in_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal2~0 (
	.dataa(curr_blk_s_1),
	.datab(\in_cnt[1]~q ),
	.datac(curr_blk_s_0),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h6996;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal2~1 (
	.dataa(Add0),
	.datab(\Equal2~0_combout ),
	.datac(Add01),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'hDFFD;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~2 (
	.dataa(\in_cnt[0]~q ),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_cnt~2_combout ),
	.cout());
defparam \in_cnt~2 .lut_mask = 16'h7777;
defparam \in_cnt~2 .sum_lutc_input = "datac";

dffeas \in_cnt[0] (
	.clk(clk),
	.d(\in_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data_p~0_combout ),
	.q(\in_cnt[0]~q ),
	.prn(vcc));
defparam \in_cnt[0] .is_wysiwyg = "true";
defparam \in_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \in_cnt~0 (
	.dataa(\in_cnt[2]~q ),
	.datab(\in_cnt[0]~q ),
	.datac(\in_cnt[1]~q ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~0_combout ),
	.cout());
defparam \in_cnt~0 .lut_mask = 16'h96FF;
defparam \in_cnt~0 .sum_lutc_input = "datac";

dffeas \in_cnt[2] (
	.clk(clk),
	.d(\in_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_data_p~0_combout ),
	.q(\in_cnt[2]~q ),
	.prn(vcc));
defparam \in_cnt[2] .is_wysiwyg = "true";
defparam \in_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \missing_sop_p~0 (
	.dataa(sink_valid),
	.datab(sink_sop),
	.datac(\in_cnt[2]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\missing_sop_p~0_combout ),
	.cout());
defparam \missing_sop_p~0 .lut_mask = 16'hBFFF;
defparam \missing_sop_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \missing_sop_p~1 (
	.dataa(\missing_sop_p~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\missing_sop_p~1_combout ),
	.cout());
defparam \missing_sop_p~1 .lut_mask = 16'hAAFF;
defparam \missing_sop_p~1 .sum_lutc_input = "datac";

dffeas missing_sop(
	.clk(clk),
	.d(\missing_sop_p~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\missing_sop~q ),
	.prn(vcc));
defparam missing_sop.is_wysiwyg = "true";
defparam missing_sop.power_up = "low";

cycloneiv_lcell_comb \unexpected_eop_p~0 (
	.dataa(sink_valid),
	.datab(sink_eop),
	.datac(gnd),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\unexpected_eop_p~0_combout ),
	.cout());
defparam \unexpected_eop_p~0 .lut_mask = 16'hEEFF;
defparam \unexpected_eop_p~0 .sum_lutc_input = "datac";

dffeas unexpected_eop(
	.clk(clk),
	.d(\unexpected_eop_p~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\unexpected_eop~q ),
	.prn(vcc));
defparam unexpected_eop.is_wysiwyg = "true";
defparam unexpected_eop.power_up = "low";

cycloneiv_lcell_comb \missing_eop_p~0 (
	.dataa(sink_valid),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(sink_eop),
	.cin(gnd),
	.combout(\missing_eop_p~0_combout ),
	.cout());
defparam \missing_eop_p~0 .lut_mask = 16'hEEFF;
defparam \missing_eop_p~0 .sum_lutc_input = "datac";

dffeas missing_eop(
	.clk(clk),
	.d(\missing_eop_p~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\missing_eop~q ),
	.prn(vcc));
defparam missing_eop.is_wysiwyg = "true";
defparam missing_eop.power_up = "low";

cycloneiv_lcell_comb \out_error_s~0 (
	.dataa(\missing_sop~q ),
	.datab(sink_error_0),
	.datac(\unexpected_eop~q ),
	.datad(\missing_eop~q ),
	.cin(gnd),
	.combout(\out_error_s~0_combout ),
	.cout());
defparam \out_error_s~0 .lut_mask = 16'hFAFC;
defparam \out_error_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_error_s~1 (
	.dataa(sink_error_1),
	.datab(\missing_eop~q ),
	.datac(\unexpected_eop~q ),
	.datad(\missing_sop~q ),
	.cin(gnd),
	.combout(\out_error_s~1_combout ),
	.cout());
defparam \out_error_s~1 .lut_mask = 16'hFAFC;
defparam \out_error_s~1 .sum_lutc_input = "datac";

dffeas \blk_shunt[2] (
	.clk(clk),
	.d(in_blk[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\blk_shunt[2]~q ),
	.prn(vcc));
defparam \blk_shunt[2] .is_wysiwyg = "true";
defparam \blk_shunt[2] .power_up = "low";

cycloneiv_lcell_comb \curr_blk_p~0 (
	.dataa(sink_sop),
	.datab(\out_data_p~0_combout ),
	.datac(gnd),
	.datad(\shunt_control~1_combout ),
	.cin(gnd),
	.combout(\curr_blk_p~0_combout ),
	.cout());
defparam \curr_blk_p~0 .lut_mask = 16'hEEFF;
defparam \curr_blk_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \curr_blk_s~2 (
	.dataa(in_blk[2]),
	.datab(\blk_shunt[2]~q ),
	.datac(gnd),
	.datad(\curr_blk_p~0_combout ),
	.cin(gnd),
	.combout(\curr_blk_s~2_combout ),
	.cout());
defparam \curr_blk_s~2 .lut_mask = 16'hAACC;
defparam \curr_blk_s~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \curr_blk_s[2]~7 (
	.dataa(sink_valid),
	.datab(\state~q ),
	.datac(source_stall_s),
	.datad(sink_sop),
	.cin(gnd),
	.combout(\curr_blk_s[2]~7_combout ),
	.cout());
defparam \curr_blk_s[2]~7 .lut_mask = 16'hFFBF;
defparam \curr_blk_s[2]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \curr_blk_s[2]~3 (
	.dataa(\state~q ),
	.datab(processing_to_end),
	.datac(\shunt_control~1_combout ),
	.datad(\curr_blk_s[2]~7_combout ),
	.cin(gnd),
	.combout(\curr_blk_s[2]~3_combout ),
	.cout());
defparam \curr_blk_s[2]~3 .lut_mask = 16'hFFBF;
defparam \curr_blk_s[2]~3 .sum_lutc_input = "datac";

dffeas \blk_shunt[1] (
	.clk(clk),
	.d(in_blk[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\blk_shunt[1]~q ),
	.prn(vcc));
defparam \blk_shunt[1] .is_wysiwyg = "true";
defparam \blk_shunt[1] .power_up = "low";

cycloneiv_lcell_comb \curr_blk_s~4 (
	.dataa(in_blk[1]),
	.datab(\blk_shunt[1]~q ),
	.datac(gnd),
	.datad(\curr_blk_p~0_combout ),
	.cin(gnd),
	.combout(\curr_blk_s~4_combout ),
	.cout());
defparam \curr_blk_s~4 .lut_mask = 16'hAACC;
defparam \curr_blk_s~4 .sum_lutc_input = "datac";

dffeas \blk_shunt[0] (
	.clk(clk),
	.d(in_blk[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\blk_shunt[0]~q ),
	.prn(vcc));
defparam \blk_shunt[0] .is_wysiwyg = "true";
defparam \blk_shunt[0] .power_up = "low";

cycloneiv_lcell_comb \curr_blk_s~5 (
	.dataa(in_blk[0]),
	.datab(\blk_shunt[0]~q ),
	.datac(gnd),
	.datad(\curr_blk_p~0_combout ),
	.cin(gnd),
	.combout(\curr_blk_s~5_combout ),
	.cout());
defparam \curr_blk_s~5 .lut_mask = 16'hAACC;
defparam \curr_blk_s~5 .sum_lutc_input = "datac";

dffeas \blk_shunt[3] (
	.clk(clk),
	.d(in_blk[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\blk_shunt[3]~q ),
	.prn(vcc));
defparam \blk_shunt[3] .is_wysiwyg = "true";
defparam \blk_shunt[3] .power_up = "low";

cycloneiv_lcell_comb \curr_blk_s~6 (
	.dataa(in_blk[3]),
	.datab(\blk_shunt[3]~q ),
	.datac(gnd),
	.datad(\curr_blk_p~0_combout ),
	.cin(gnd),
	.combout(\curr_blk_s~6_combout ),
	.cout());
defparam \curr_blk_s~6 .lut_mask = 16'hAACC;
defparam \curr_blk_s~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb in_pwr_2(
	.dataa(in_blk[1]),
	.datab(in_blk[3]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_pwr_2~combout ),
	.cout());
defparam in_pwr_2.lut_mask = 16'hEEEE;
defparam in_pwr_2.sum_lutc_input = "datac";

dffeas pwr_2_shunt(
	.clk(clk),
	.d(\in_pwr_2~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\pwr_2_shunt~q ),
	.prn(vcc));
defparam pwr_2_shunt.is_wysiwyg = "true";
defparam pwr_2_shunt.power_up = "low";

cycloneiv_lcell_comb \curr_pwr_2_s~0 (
	.dataa(\pwr_2_shunt~q ),
	.datab(\curr_blk_p~0_combout ),
	.datac(in_blk[1]),
	.datad(in_blk[3]),
	.cin(gnd),
	.combout(\curr_pwr_2_s~0_combout ),
	.cout());
defparam \curr_pwr_2_s~0 .lut_mask = 16'hFFB8;
defparam \curr_pwr_2_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \leaving_s5_state~0 (
	.dataa(\state~q ),
	.datab(gnd),
	.datac(source_stall_s),
	.datad(processing_to_end),
	.cin(gnd),
	.combout(\leaving_s5_state~0_combout ),
	.cout());
defparam \leaving_s5_state~0 .lut_mask = 16'hAFFF;
defparam \leaving_s5_state~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_valid_s~0 (
	.dataa(\leaving_s5_state~0_combout ),
	.datab(\out_data_p~0_combout ),
	.datac(gnd),
	.datad(\shunt_control~1_combout ),
	.cin(gnd),
	.combout(\out_valid_s~0_combout ),
	.cout());
defparam \out_valid_s~0 .lut_mask = 16'hEEFF;
defparam \out_valid_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \got_sop~0 (
	.dataa(\got_sop~q ),
	.datab(sink_sop),
	.datac(\out_data_p~0_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\got_sop~0_combout ),
	.cout());
defparam \got_sop~0 .lut_mask = 16'hACFF;
defparam \got_sop~0 .sum_lutc_input = "datac";

dffeas got_sop(
	.clk(clk),
	.d(\got_sop~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\got_sop~q ),
	.prn(vcc));
defparam got_sop.is_wysiwyg = "true";
defparam got_sop.power_up = "low";

cycloneiv_lcell_comb \out_valid_s~1 (
	.dataa(\out_valid_s~0_combout ),
	.datab(sink_sop),
	.datac(\got_sop~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_s~1_combout ),
	.cout());
defparam \out_valid_s~1 .lut_mask = 16'hFEFE;
defparam \out_valid_s~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt~0 (
	.dataa(gnd),
	.datab(cnt_0),
	.datac(cnt_1),
	.datad(Equal1),
	.cin(gnd),
	.combout(\cnt~0_combout ),
	.cout());
defparam \cnt~0 .lut_mask = 16'hFF3C;
defparam \cnt~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt~1 (
	.dataa(cnt_0),
	.datab(Equal1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\cnt~1_combout ),
	.cout());
defparam \cnt~1 .lut_mask = 16'hDDDD;
defparam \cnt~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt~2 (
	.dataa(cnt_2),
	.datab(cnt_0),
	.datac(cnt_1),
	.datad(Equal1),
	.cin(gnd),
	.combout(\cnt~2_combout ),
	.cout());
defparam \cnt~2 .lut_mask = 16'hFF96;
defparam \cnt~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal1~0 (
	.dataa(curr_blk_s_1),
	.datab(cnt_1),
	.datac(curr_blk_s_0),
	.datad(cnt_0),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h6996;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \entering_s5_state~1 (
	.dataa(entering_s5_state),
	.datab(\shunt_control~0_combout ),
	.datac(\Equal5~0_combout ),
	.datad(\Equal5~1_combout ),
	.cin(gnd),
	.combout(\entering_s5_state~1_combout ),
	.cout());
defparam \entering_s5_state~1 .lut_mask = 16'hEFFF;
defparam \entering_s5_state~1 .sum_lutc_input = "datac";

dffeas \in_data_shunt[8] (
	.clk(clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[8]~q ),
	.prn(vcc));
defparam \in_data_shunt[8] .is_wysiwyg = "true";
defparam \in_data_shunt[8] .power_up = "low";

cycloneiv_lcell_comb \out_data~0 (
	.dataa(\in_data_shunt[8]~q ),
	.datab(in_data[8]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~0_combout ),
	.cout());
defparam \out_data~0 .lut_mask = 16'hAACC;
defparam \out_data~0 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[0]~q ),
	.prn(vcc));
defparam \in_data_shunt[0] .is_wysiwyg = "true";
defparam \in_data_shunt[0] .power_up = "low";

cycloneiv_lcell_comb \out_data~1 (
	.dataa(\in_data_shunt[0]~q ),
	.datab(in_data[0]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~1_combout ),
	.cout());
defparam \out_data~1 .lut_mask = 16'hAACC;
defparam \out_data~1 .sum_lutc_input = "datac";

dffeas inverse_shunt(
	.clk(clk),
	.d(in_inverse),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\inverse_shunt~q ),
	.prn(vcc));
defparam inverse_shunt.is_wysiwyg = "true";
defparam inverse_shunt.power_up = "low";

cycloneiv_lcell_comb \curr_inverse_s~0 (
	.dataa(in_inverse),
	.datab(\inverse_shunt~q ),
	.datac(gnd),
	.datad(\curr_blk_p~0_combout ),
	.cin(gnd),
	.combout(\curr_inverse_s~0_combout ),
	.cout());
defparam \curr_inverse_s~0 .lut_mask = 16'hAACC;
defparam \curr_inverse_s~0 .sum_lutc_input = "datac";

dffeas \in_data_shunt[9] (
	.clk(clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[9]~q ),
	.prn(vcc));
defparam \in_data_shunt[9] .is_wysiwyg = "true";
defparam \in_data_shunt[9] .power_up = "low";

cycloneiv_lcell_comb \out_data~2 (
	.dataa(\in_data_shunt[9]~q ),
	.datab(in_data[9]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~2_combout ),
	.cout());
defparam \out_data~2 .lut_mask = 16'hAACC;
defparam \out_data~2 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[1]~q ),
	.prn(vcc));
defparam \in_data_shunt[1] .is_wysiwyg = "true";
defparam \in_data_shunt[1] .power_up = "low";

cycloneiv_lcell_comb \out_data~3 (
	.dataa(\in_data_shunt[1]~q ),
	.datab(in_data[1]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~3_combout ),
	.cout());
defparam \out_data~3 .lut_mask = 16'hAACC;
defparam \out_data~3 .sum_lutc_input = "datac";

dffeas \in_data_shunt[10] (
	.clk(clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[10]~q ),
	.prn(vcc));
defparam \in_data_shunt[10] .is_wysiwyg = "true";
defparam \in_data_shunt[10] .power_up = "low";

cycloneiv_lcell_comb \out_data~4 (
	.dataa(\in_data_shunt[10]~q ),
	.datab(in_data[10]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~4_combout ),
	.cout());
defparam \out_data~4 .lut_mask = 16'hAACC;
defparam \out_data~4 .sum_lutc_input = "datac";

dffeas \in_data_shunt[2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[2]~q ),
	.prn(vcc));
defparam \in_data_shunt[2] .is_wysiwyg = "true";
defparam \in_data_shunt[2] .power_up = "low";

cycloneiv_lcell_comb \out_data~5 (
	.dataa(\in_data_shunt[2]~q ),
	.datab(in_data[2]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~5_combout ),
	.cout());
defparam \out_data~5 .lut_mask = 16'hAACC;
defparam \out_data~5 .sum_lutc_input = "datac";

dffeas \in_data_shunt[11] (
	.clk(clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[11]~q ),
	.prn(vcc));
defparam \in_data_shunt[11] .is_wysiwyg = "true";
defparam \in_data_shunt[11] .power_up = "low";

cycloneiv_lcell_comb \out_data~6 (
	.dataa(\in_data_shunt[11]~q ),
	.datab(in_data[11]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~6_combout ),
	.cout());
defparam \out_data~6 .lut_mask = 16'hAACC;
defparam \out_data~6 .sum_lutc_input = "datac";

dffeas \in_data_shunt[3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[3]~q ),
	.prn(vcc));
defparam \in_data_shunt[3] .is_wysiwyg = "true";
defparam \in_data_shunt[3] .power_up = "low";

cycloneiv_lcell_comb \out_data~7 (
	.dataa(\in_data_shunt[3]~q ),
	.datab(in_data[3]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~7_combout ),
	.cout());
defparam \out_data~7 .lut_mask = 16'hAACC;
defparam \out_data~7 .sum_lutc_input = "datac";

dffeas \in_data_shunt[12] (
	.clk(clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[12]~q ),
	.prn(vcc));
defparam \in_data_shunt[12] .is_wysiwyg = "true";
defparam \in_data_shunt[12] .power_up = "low";

cycloneiv_lcell_comb \out_data~8 (
	.dataa(\in_data_shunt[12]~q ),
	.datab(in_data[12]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~8_combout ),
	.cout());
defparam \out_data~8 .lut_mask = 16'hAACC;
defparam \out_data~8 .sum_lutc_input = "datac";

dffeas \in_data_shunt[4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[4]~q ),
	.prn(vcc));
defparam \in_data_shunt[4] .is_wysiwyg = "true";
defparam \in_data_shunt[4] .power_up = "low";

cycloneiv_lcell_comb \out_data~9 (
	.dataa(\in_data_shunt[4]~q ),
	.datab(in_data[4]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~9_combout ),
	.cout());
defparam \out_data~9 .lut_mask = 16'hAACC;
defparam \out_data~9 .sum_lutc_input = "datac";

dffeas \in_data_shunt[13] (
	.clk(clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[13]~q ),
	.prn(vcc));
defparam \in_data_shunt[13] .is_wysiwyg = "true";
defparam \in_data_shunt[13] .power_up = "low";

cycloneiv_lcell_comb \out_data~10 (
	.dataa(\in_data_shunt[13]~q ),
	.datab(in_data[13]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~10_combout ),
	.cout());
defparam \out_data~10 .lut_mask = 16'hAACC;
defparam \out_data~10 .sum_lutc_input = "datac";

dffeas \in_data_shunt[5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[5]~q ),
	.prn(vcc));
defparam \in_data_shunt[5] .is_wysiwyg = "true";
defparam \in_data_shunt[5] .power_up = "low";

cycloneiv_lcell_comb \out_data~11 (
	.dataa(\in_data_shunt[5]~q ),
	.datab(in_data[5]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~11_combout ),
	.cout());
defparam \out_data~11 .lut_mask = 16'hAACC;
defparam \out_data~11 .sum_lutc_input = "datac";

dffeas \in_data_shunt[14] (
	.clk(clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[14]~q ),
	.prn(vcc));
defparam \in_data_shunt[14] .is_wysiwyg = "true";
defparam \in_data_shunt[14] .power_up = "low";

cycloneiv_lcell_comb \out_data~12 (
	.dataa(\in_data_shunt[14]~q ),
	.datab(in_data[14]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~12_combout ),
	.cout());
defparam \out_data~12 .lut_mask = 16'hAACC;
defparam \out_data~12 .sum_lutc_input = "datac";

dffeas \in_data_shunt[6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[6]~q ),
	.prn(vcc));
defparam \in_data_shunt[6] .is_wysiwyg = "true";
defparam \in_data_shunt[6] .power_up = "low";

cycloneiv_lcell_comb \out_data~13 (
	.dataa(\in_data_shunt[6]~q ),
	.datab(in_data[6]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~13_combout ),
	.cout());
defparam \out_data~13 .lut_mask = 16'hAACC;
defparam \out_data~13 .sum_lutc_input = "datac";

dffeas \in_data_shunt[15] (
	.clk(clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[15]~q ),
	.prn(vcc));
defparam \in_data_shunt[15] .is_wysiwyg = "true";
defparam \in_data_shunt[15] .power_up = "low";

cycloneiv_lcell_comb \out_data~14 (
	.dataa(\in_data_shunt[15]~q ),
	.datab(in_data[15]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~14_combout ),
	.cout());
defparam \out_data~14 .lut_mask = 16'hAACC;
defparam \out_data~14 .sum_lutc_input = "datac";

dffeas \in_data_shunt[7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\entering_s5_state~1_combout ),
	.q(\in_data_shunt[7]~q ),
	.prn(vcc));
defparam \in_data_shunt[7] .is_wysiwyg = "true";
defparam \in_data_shunt[7] .power_up = "low";

cycloneiv_lcell_comb \out_data~15 (
	.dataa(\in_data_shunt[7]~q ),
	.datab(in_data[7]),
	.datac(gnd),
	.datad(\leaving_s5_state~0_combout ),
	.cin(gnd),
	.combout(\out_data~15_combout ),
	.cout());
defparam \out_data~15 .lut_mask = 16'hAACC;
defparam \out_data~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_input_sel[0]~0 (
	.dataa(in_blk[2]),
	.datab(in_blk[3]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_input_sel[0]~0_combout ),
	.cout());
defparam \stg_input_sel[0]~0 .lut_mask = 16'hEEEE;
defparam \stg_input_sel[0]~0 .sum_lutc_input = "datac";

dffeas \input_sel_shunt[0] (
	.clk(clk),
	.d(\stg_input_sel[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_control~1_combout ),
	.q(\input_sel_shunt[0]~q ),
	.prn(vcc));
defparam \input_sel_shunt[0] .is_wysiwyg = "true";
defparam \input_sel_shunt[0] .power_up = "low";

cycloneiv_lcell_comb \curr_input_sel_s~0 (
	.dataa(\input_sel_shunt[0]~q ),
	.datab(\curr_blk_p~0_combout ),
	.datac(in_blk[2]),
	.datad(in_blk[3]),
	.cin(gnd),
	.combout(\curr_input_sel_s~0_combout ),
	.cout());
defparam \curr_input_sel_s~0 .lut_mask = 16'hFFB8;
defparam \curr_input_sel_s~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_avalon_streaming_block_source (
	in_data,
	source_stall_s1,
	stateIDLE,
	Equal0,
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Add0,
	Add01,
	Equal1,
	source_data_0,
	source_data_1,
	source_data_2,
	source_data_3,
	source_data_4,
	source_data_5,
	source_data_6,
	source_data_7,
	source_data_8,
	source_data_9,
	source_data_10,
	source_data_11,
	source_data_12,
	source_data_13,
	source_data_14,
	source_data_15,
	rd_valid_dd,
	rd_enable,
	out_valid,
	out_enable,
	stall_p,
	Add02,
	out_valid1,
	out_valid2,
	clk,
	reset,
	source_ready)/* synthesis synthesis_greybox=1 */;
input 	[15:0] in_data;
output 	source_stall_s1;
output 	stateIDLE;
output 	Equal0;
input 	curr_blk_s_2;
input 	curr_blk_s_1;
input 	curr_blk_s_0;
input 	curr_blk_s_3;
output 	Add0;
output 	Add01;
output 	Equal1;
output 	source_data_0;
output 	source_data_1;
output 	source_data_2;
output 	source_data_3;
output 	source_data_4;
output 	source_data_5;
output 	source_data_6;
output 	source_data_7;
output 	source_data_8;
output 	source_data_9;
output 	source_data_10;
output 	source_data_11;
output 	source_data_12;
output 	source_data_13;
output 	source_data_14;
output 	source_data_15;
input 	rd_valid_dd;
input 	rd_enable;
input 	out_valid;
input 	out_enable;
output 	stall_p;
output 	Add02;
input 	out_valid1;
input 	out_valid2;
input 	clk;
input 	reset;
input 	source_ready;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \Selector1~0_combout ;
wire \Selector1~1_combout ;
wire \state.OUT_1~q ;
wire \Selector2~0_combout ;
wire \Selector2~1_combout ;
wire \state.OUT_2~q ;
wire \Selector3~0_combout ;
wire \state.OUT_3~q ;
wire \stall_p~1_combout ;
wire \out_data_p~0_combout ;
wire \Selector0~0_combout ;
wire \data_count~0_combout ;
wire \data_count[0]~q ;
wire \data_count~3_combout ;
wire \data_count[1]~q ;
wire \data_count~2_combout ;
wire \data_count[2]~q ;
wire \Add1~0_combout ;
wire \data_count~1_combout ;
wire \data_count[3]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \shunt_p~2_combout ;
wire \in_data_shunt[1][0]~q ;
wire \shunt_p~0_combout ;
wire \shunt_p~1_combout ;
wire \in_data_shunt~0_combout ;
wire \in_data_shunt[0][4]~1_combout ;
wire \in_data_shunt[0][4]~2_combout ;
wire \in_data_shunt[0][0]~q ;
wire \out_data_p~1_combout ;
wire \source_data~0_combout ;
wire \source_data[6]~1_combout ;
wire \source_data[6]~2_combout ;
wire \in_data_shunt[1][1]~q ;
wire \in_data_shunt~3_combout ;
wire \in_data_shunt[0][1]~q ;
wire \source_data~3_combout ;
wire \in_data_shunt[1][2]~q ;
wire \in_data_shunt~4_combout ;
wire \in_data_shunt[0][2]~q ;
wire \source_data~4_combout ;
wire \in_data_shunt[1][3]~q ;
wire \in_data_shunt~5_combout ;
wire \in_data_shunt[0][3]~q ;
wire \source_data~5_combout ;
wire \in_data_shunt[1][4]~q ;
wire \in_data_shunt~6_combout ;
wire \in_data_shunt[0][4]~q ;
wire \source_data~6_combout ;
wire \in_data_shunt[1][5]~q ;
wire \in_data_shunt~7_combout ;
wire \in_data_shunt[0][5]~q ;
wire \source_data~7_combout ;
wire \in_data_shunt[1][6]~q ;
wire \in_data_shunt~8_combout ;
wire \in_data_shunt[0][6]~q ;
wire \source_data~8_combout ;
wire \in_data_shunt[1][7]~q ;
wire \in_data_shunt~9_combout ;
wire \in_data_shunt[0][7]~q ;
wire \source_data~9_combout ;
wire \in_data_shunt[1][8]~q ;
wire \in_data_shunt~10_combout ;
wire \in_data_shunt[0][8]~q ;
wire \source_data~10_combout ;
wire \in_data_shunt[1][9]~q ;
wire \in_data_shunt~11_combout ;
wire \in_data_shunt[0][9]~q ;
wire \source_data~11_combout ;
wire \in_data_shunt[1][10]~q ;
wire \in_data_shunt~12_combout ;
wire \in_data_shunt[0][10]~q ;
wire \source_data~12_combout ;
wire \in_data_shunt[1][11]~q ;
wire \in_data_shunt~13_combout ;
wire \in_data_shunt[0][11]~q ;
wire \source_data~13_combout ;
wire \in_data_shunt[1][12]~q ;
wire \in_data_shunt~14_combout ;
wire \in_data_shunt[0][12]~q ;
wire \source_data~14_combout ;
wire \in_data_shunt[1][13]~q ;
wire \in_data_shunt~15_combout ;
wire \in_data_shunt[0][13]~q ;
wire \source_data~15_combout ;
wire \in_data_shunt[1][14]~q ;
wire \in_data_shunt~16_combout ;
wire \in_data_shunt[0][14]~q ;
wire \source_data~16_combout ;
wire \in_data_shunt[1][15]~q ;
wire \in_data_shunt~17_combout ;
wire \in_data_shunt[0][15]~q ;
wire \source_data~17_combout ;


dffeas source_stall_s(
	.clk(clk),
	.d(\stall_p~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(source_stall_s1),
	.prn(vcc));
defparam source_stall_s.is_wysiwyg = "true";
defparam source_stall_s.power_up = "low";

dffeas \state.IDLE (
	.clk(clk),
	.d(\Selector0~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(stateIDLE),
	.prn(vcc));
defparam \state.IDLE .is_wysiwyg = "true";
defparam \state.IDLE .power_up = "low";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(\data_count[0]~q ),
	.datab(\data_count[3]~q ),
	.datac(\data_count[2]~q ),
	.datad(\data_count[1]~q ),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h7FFF;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~0 (
	.dataa(curr_blk_s_2),
	.datab(curr_blk_s_1),
	.datac(curr_blk_s_0),
	.datad(curr_blk_s_3),
	.cin(gnd),
	.combout(Add0),
	.cout());
defparam \Add0~0 .lut_mask = 16'h6996;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~1 (
	.dataa(gnd),
	.datab(curr_blk_s_1),
	.datac(curr_blk_s_0),
	.datad(curr_blk_s_2),
	.cin(gnd),
	.combout(Add01),
	.cout());
defparam \Add0~1 .lut_mask = 16'hC33C;
defparam \Add0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal1~2 (
	.dataa(\Equal1~0_combout ),
	.datab(\Equal1~1_combout ),
	.datac(\data_count[2]~q ),
	.datad(Add01),
	.cin(gnd),
	.combout(Equal1),
	.cout());
defparam \Equal1~2 .lut_mask = 16'hEFFE;
defparam \Equal1~2 .sum_lutc_input = "datac";

dffeas \source_data[0] (
	.clk(clk),
	.d(\source_data~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_0),
	.prn(vcc));
defparam \source_data[0] .is_wysiwyg = "true";
defparam \source_data[0] .power_up = "low";

dffeas \source_data[1] (
	.clk(clk),
	.d(\source_data~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_1),
	.prn(vcc));
defparam \source_data[1] .is_wysiwyg = "true";
defparam \source_data[1] .power_up = "low";

dffeas \source_data[2] (
	.clk(clk),
	.d(\source_data~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_2),
	.prn(vcc));
defparam \source_data[2] .is_wysiwyg = "true";
defparam \source_data[2] .power_up = "low";

dffeas \source_data[3] (
	.clk(clk),
	.d(\source_data~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_3),
	.prn(vcc));
defparam \source_data[3] .is_wysiwyg = "true";
defparam \source_data[3] .power_up = "low";

dffeas \source_data[4] (
	.clk(clk),
	.d(\source_data~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_4),
	.prn(vcc));
defparam \source_data[4] .is_wysiwyg = "true";
defparam \source_data[4] .power_up = "low";

dffeas \source_data[5] (
	.clk(clk),
	.d(\source_data~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_5),
	.prn(vcc));
defparam \source_data[5] .is_wysiwyg = "true";
defparam \source_data[5] .power_up = "low";

dffeas \source_data[6] (
	.clk(clk),
	.d(\source_data~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_6),
	.prn(vcc));
defparam \source_data[6] .is_wysiwyg = "true";
defparam \source_data[6] .power_up = "low";

dffeas \source_data[7] (
	.clk(clk),
	.d(\source_data~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_7),
	.prn(vcc));
defparam \source_data[7] .is_wysiwyg = "true";
defparam \source_data[7] .power_up = "low";

dffeas \source_data[8] (
	.clk(clk),
	.d(\source_data~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_8),
	.prn(vcc));
defparam \source_data[8] .is_wysiwyg = "true";
defparam \source_data[8] .power_up = "low";

dffeas \source_data[9] (
	.clk(clk),
	.d(\source_data~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_9),
	.prn(vcc));
defparam \source_data[9] .is_wysiwyg = "true";
defparam \source_data[9] .power_up = "low";

dffeas \source_data[10] (
	.clk(clk),
	.d(\source_data~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_10),
	.prn(vcc));
defparam \source_data[10] .is_wysiwyg = "true";
defparam \source_data[10] .power_up = "low";

dffeas \source_data[11] (
	.clk(clk),
	.d(\source_data~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_11),
	.prn(vcc));
defparam \source_data[11] .is_wysiwyg = "true";
defparam \source_data[11] .power_up = "low";

dffeas \source_data[12] (
	.clk(clk),
	.d(\source_data~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_12),
	.prn(vcc));
defparam \source_data[12] .is_wysiwyg = "true";
defparam \source_data[12] .power_up = "low";

dffeas \source_data[13] (
	.clk(clk),
	.d(\source_data~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_13),
	.prn(vcc));
defparam \source_data[13] .is_wysiwyg = "true";
defparam \source_data[13] .power_up = "low";

dffeas \source_data[14] (
	.clk(clk),
	.d(\source_data~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_14),
	.prn(vcc));
defparam \source_data[14] .is_wysiwyg = "true";
defparam \source_data[14] .power_up = "low";

dffeas \source_data[15] (
	.clk(clk),
	.d(\source_data~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\source_data[6]~2_combout ),
	.q(source_data_15),
	.prn(vcc));
defparam \source_data[15] .is_wysiwyg = "true";
defparam \source_data[15] .power_up = "low";

cycloneiv_lcell_comb \stall_p~2 (
	.dataa(stateIDLE),
	.datab(source_ready),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(stall_p),
	.cout());
defparam \stall_p~2 .lut_mask = 16'hEEEE;
defparam \stall_p~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(curr_blk_s_1),
	.datad(curr_blk_s_0),
	.cin(gnd),
	.combout(Add02),
	.cout());
defparam \Add0~2 .lut_mask = 16'h0FF0;
defparam \Add0~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Selector1~0 (
	.dataa(source_ready),
	.datab(\state.OUT_2~q ),
	.datac(out_valid2),
	.datad(stateIDLE),
	.cin(gnd),
	.combout(\Selector1~0_combout ),
	.cout());
defparam \Selector1~0 .lut_mask = 16'hACFF;
defparam \Selector1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Selector1~1 (
	.dataa(\Selector1~0_combout ),
	.datab(\state.OUT_1~q ),
	.datac(source_ready),
	.datad(out_valid2),
	.cin(gnd),
	.combout(\Selector1~1_combout ),
	.cout());
defparam \Selector1~1 .lut_mask = 16'hEFFE;
defparam \Selector1~1 .sum_lutc_input = "datac";

dffeas \state.OUT_1 (
	.clk(clk),
	.d(\Selector1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.OUT_1~q ),
	.prn(vcc));
defparam \state.OUT_1 .is_wysiwyg = "true";
defparam \state.OUT_1 .power_up = "low";

cycloneiv_lcell_comb \Selector2~0 (
	.dataa(source_ready),
	.datab(\state.OUT_1~q ),
	.datac(\state.OUT_3~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Selector2~0_combout ),
	.cout());
defparam \Selector2~0 .lut_mask = 16'hD8D8;
defparam \Selector2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Selector2~1 (
	.dataa(\state.OUT_2~q ),
	.datab(source_ready),
	.datac(out_valid2),
	.datad(\Selector2~0_combout ),
	.cin(gnd),
	.combout(\Selector2~1_combout ),
	.cout());
defparam \Selector2~1 .lut_mask = 16'hFFBE;
defparam \Selector2~1 .sum_lutc_input = "datac";

dffeas \state.OUT_2 (
	.clk(clk),
	.d(\Selector2~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.OUT_2~q ),
	.prn(vcc));
defparam \state.OUT_2 .is_wysiwyg = "true";
defparam \state.OUT_2 .power_up = "low";

cycloneiv_lcell_comb \Selector3~0 (
	.dataa(\state.OUT_3~q ),
	.datab(out_valid2),
	.datac(\state.OUT_2~q ),
	.datad(source_ready),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
defparam \Selector3~0 .lut_mask = 16'hFEFF;
defparam \Selector3~0 .sum_lutc_input = "datac";

dffeas \state.OUT_3 (
	.clk(clk),
	.d(\Selector3~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\state.OUT_3~q ),
	.prn(vcc));
defparam \state.OUT_3 .is_wysiwyg = "true";
defparam \state.OUT_3 .power_up = "low";

cycloneiv_lcell_comb \stall_p~1 (
	.dataa(stateIDLE),
	.datab(\state.OUT_3~q ),
	.datac(gnd),
	.datad(source_ready),
	.cin(gnd),
	.combout(\stall_p~1_combout ),
	.cout());
defparam \stall_p~1 .lut_mask = 16'hEEFF;
defparam \stall_p~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_data_p~0 (
	.dataa(source_ready),
	.datab(\state.OUT_1~q ),
	.datac(gnd),
	.datad(stateIDLE),
	.cin(gnd),
	.combout(\out_data_p~0_combout ),
	.cout());
defparam \out_data_p~0 .lut_mask = 16'hEEFF;
defparam \out_data_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Selector0~0 (
	.dataa(\out_data_p~0_combout ),
	.datab(gnd),
	.datac(rd_valid_dd),
	.datad(out_valid1),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
defparam \Selector0~0 .lut_mask = 16'hFFF5;
defparam \Selector0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \data_count~0 (
	.dataa(\data_count[0]~q ),
	.datab(Equal1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\data_count~0_combout ),
	.cout());
defparam \data_count~0 .lut_mask = 16'h7777;
defparam \data_count~0 .sum_lutc_input = "datac";

dffeas \data_count[0] (
	.clk(clk),
	.d(\data_count~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(stall_p),
	.q(\data_count[0]~q ),
	.prn(vcc));
defparam \data_count[0] .is_wysiwyg = "true";
defparam \data_count[0] .power_up = "low";

cycloneiv_lcell_comb \data_count~3 (
	.dataa(gnd),
	.datab(\data_count[0]~q ),
	.datac(\data_count[1]~q ),
	.datad(Equal1),
	.cin(gnd),
	.combout(\data_count~3_combout ),
	.cout());
defparam \data_count~3 .lut_mask = 16'h3CFF;
defparam \data_count~3 .sum_lutc_input = "datac";

dffeas \data_count[1] (
	.clk(clk),
	.d(\data_count~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(stall_p),
	.q(\data_count[1]~q ),
	.prn(vcc));
defparam \data_count[1] .is_wysiwyg = "true";
defparam \data_count[1] .power_up = "low";

cycloneiv_lcell_comb \data_count~2 (
	.dataa(\data_count[2]~q ),
	.datab(\data_count[0]~q ),
	.datac(\data_count[1]~q ),
	.datad(Equal1),
	.cin(gnd),
	.combout(\data_count~2_combout ),
	.cout());
defparam \data_count~2 .lut_mask = 16'h96FF;
defparam \data_count~2 .sum_lutc_input = "datac";

dffeas \data_count[2] (
	.clk(clk),
	.d(\data_count~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(stall_p),
	.q(\data_count[2]~q ),
	.prn(vcc));
defparam \data_count[2] .is_wysiwyg = "true";
defparam \data_count[2] .power_up = "low";

cycloneiv_lcell_comb \Add1~0 (
	.dataa(\data_count[3]~q ),
	.datab(\data_count[0]~q ),
	.datac(\data_count[2]~q ),
	.datad(\data_count[1]~q ),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6996;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \data_count~1 (
	.dataa(\Add1~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(Equal1),
	.cin(gnd),
	.combout(\data_count~1_combout ),
	.cout());
defparam \data_count~1 .lut_mask = 16'hAAFF;
defparam \data_count~1 .sum_lutc_input = "datac";

dffeas \data_count[3] (
	.clk(clk),
	.d(\data_count~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(stall_p),
	.q(\data_count[3]~q ),
	.prn(vcc));
defparam \data_count[3] .is_wysiwyg = "true";
defparam \data_count[3] .power_up = "low";

cycloneiv_lcell_comb \Equal1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\data_count[3]~q ),
	.datad(Add0),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h0FF0;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal1~1 (
	.dataa(\data_count[1]~q ),
	.datab(curr_blk_s_1),
	.datac(curr_blk_s_0),
	.datad(\data_count[0]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'h6996;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shunt_p~2 (
	.dataa(rd_valid_dd),
	.datab(out_valid1),
	.datac(\state.OUT_2~q ),
	.datad(source_ready),
	.cin(gnd),
	.combout(\shunt_p~2_combout ),
	.cout());
defparam \shunt_p~2 .lut_mask = 16'hFEFF;
defparam \shunt_p~2 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][0] (
	.clk(clk),
	.d(in_data[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][0]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][0] .is_wysiwyg = "true";
defparam \in_data_shunt[1][0] .power_up = "low";

cycloneiv_lcell_comb \shunt_p~0 (
	.dataa(rd_valid_dd),
	.datab(\state.OUT_2~q ),
	.datac(\state.OUT_1~q ),
	.datad(source_ready),
	.cin(gnd),
	.combout(\shunt_p~0_combout ),
	.cout());
defparam \shunt_p~0 .lut_mask = 16'hFAFC;
defparam \shunt_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shunt_p~1 (
	.dataa(rd_enable),
	.datab(out_valid),
	.datac(out_enable),
	.datad(\shunt_p~0_combout ),
	.cin(gnd),
	.combout(\shunt_p~1_combout ),
	.cout());
defparam \shunt_p~1 .lut_mask = 16'hFFFE;
defparam \shunt_p~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_data_shunt~0 (
	.dataa(in_data[0]),
	.datab(\in_data_shunt[1][0]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~0_combout ),
	.cout());
defparam \in_data_shunt~0 .lut_mask = 16'hAACC;
defparam \in_data_shunt~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_data_shunt[0][4]~1 (
	.dataa(\state.OUT_2~q ),
	.datab(\state.OUT_1~q ),
	.datac(source_ready),
	.datad(rd_valid_dd),
	.cin(gnd),
	.combout(\in_data_shunt[0][4]~1_combout ),
	.cout());
defparam \in_data_shunt[0][4]~1 .lut_mask = 16'h53FF;
defparam \in_data_shunt[0][4]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_data_shunt[0][4]~2 (
	.dataa(source_ready),
	.datab(\state.OUT_3~q ),
	.datac(out_valid1),
	.datad(\in_data_shunt[0][4]~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt[0][4]~2_combout ),
	.cout());
defparam \in_data_shunt[0][4]~2 .lut_mask = 16'hFEFF;
defparam \in_data_shunt[0][4]~2 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][0] (
	.clk(clk),
	.d(\in_data_shunt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][0]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][0] .is_wysiwyg = "true";
defparam \in_data_shunt[0][0] .power_up = "low";

cycloneiv_lcell_comb \out_data_p~1 (
	.dataa(rd_valid_dd),
	.datab(out_valid1),
	.datac(\out_data_p~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_data_p~1_combout ),
	.cout());
defparam \out_data_p~1 .lut_mask = 16'hFEFE;
defparam \out_data_p~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_data~0 (
	.dataa(in_data[0]),
	.datab(\in_data_shunt[0][0]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~0_combout ),
	.cout());
defparam \source_data~0 .lut_mask = 16'hAACC;
defparam \source_data~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_data[6]~1 (
	.dataa(\state.OUT_3~q ),
	.datab(\state.OUT_2~q ),
	.datac(source_ready),
	.datad(gnd),
	.cin(gnd),
	.combout(\source_data[6]~1_combout ),
	.cout());
defparam \source_data[6]~1 .lut_mask = 16'h7F7F;
defparam \source_data[6]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \source_data[6]~2 (
	.dataa(rd_valid_dd),
	.datab(out_valid1),
	.datac(\out_data_p~0_combout ),
	.datad(\source_data[6]~1_combout ),
	.cin(gnd),
	.combout(\source_data[6]~2_combout ),
	.cout());
defparam \source_data[6]~2 .lut_mask = 16'hFEFF;
defparam \source_data[6]~2 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][1] (
	.clk(clk),
	.d(in_data[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][1]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][1] .is_wysiwyg = "true";
defparam \in_data_shunt[1][1] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~3 (
	.dataa(in_data[1]),
	.datab(\in_data_shunt[1][1]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~3_combout ),
	.cout());
defparam \in_data_shunt~3 .lut_mask = 16'hAACC;
defparam \in_data_shunt~3 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][1] (
	.clk(clk),
	.d(\in_data_shunt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][1]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][1] .is_wysiwyg = "true";
defparam \in_data_shunt[0][1] .power_up = "low";

cycloneiv_lcell_comb \source_data~3 (
	.dataa(in_data[1]),
	.datab(\in_data_shunt[0][1]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~3_combout ),
	.cout());
defparam \source_data~3 .lut_mask = 16'hAACC;
defparam \source_data~3 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][2] (
	.clk(clk),
	.d(in_data[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][2]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][2] .is_wysiwyg = "true";
defparam \in_data_shunt[1][2] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~4 (
	.dataa(in_data[2]),
	.datab(\in_data_shunt[1][2]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~4_combout ),
	.cout());
defparam \in_data_shunt~4 .lut_mask = 16'hAACC;
defparam \in_data_shunt~4 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][2] (
	.clk(clk),
	.d(\in_data_shunt~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][2]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][2] .is_wysiwyg = "true";
defparam \in_data_shunt[0][2] .power_up = "low";

cycloneiv_lcell_comb \source_data~4 (
	.dataa(in_data[2]),
	.datab(\in_data_shunt[0][2]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~4_combout ),
	.cout());
defparam \source_data~4 .lut_mask = 16'hAACC;
defparam \source_data~4 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][3] (
	.clk(clk),
	.d(in_data[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][3]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][3] .is_wysiwyg = "true";
defparam \in_data_shunt[1][3] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~5 (
	.dataa(in_data[3]),
	.datab(\in_data_shunt[1][3]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~5_combout ),
	.cout());
defparam \in_data_shunt~5 .lut_mask = 16'hAACC;
defparam \in_data_shunt~5 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][3] (
	.clk(clk),
	.d(\in_data_shunt~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][3]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][3] .is_wysiwyg = "true";
defparam \in_data_shunt[0][3] .power_up = "low";

cycloneiv_lcell_comb \source_data~5 (
	.dataa(in_data[3]),
	.datab(\in_data_shunt[0][3]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~5_combout ),
	.cout());
defparam \source_data~5 .lut_mask = 16'hAACC;
defparam \source_data~5 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][4] (
	.clk(clk),
	.d(in_data[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][4]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][4] .is_wysiwyg = "true";
defparam \in_data_shunt[1][4] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~6 (
	.dataa(in_data[4]),
	.datab(\in_data_shunt[1][4]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~6_combout ),
	.cout());
defparam \in_data_shunt~6 .lut_mask = 16'hAACC;
defparam \in_data_shunt~6 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][4] (
	.clk(clk),
	.d(\in_data_shunt~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][4]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][4] .is_wysiwyg = "true";
defparam \in_data_shunt[0][4] .power_up = "low";

cycloneiv_lcell_comb \source_data~6 (
	.dataa(in_data[4]),
	.datab(\in_data_shunt[0][4]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~6_combout ),
	.cout());
defparam \source_data~6 .lut_mask = 16'hAACC;
defparam \source_data~6 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][5] (
	.clk(clk),
	.d(in_data[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][5]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][5] .is_wysiwyg = "true";
defparam \in_data_shunt[1][5] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~7 (
	.dataa(in_data[5]),
	.datab(\in_data_shunt[1][5]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~7_combout ),
	.cout());
defparam \in_data_shunt~7 .lut_mask = 16'hAACC;
defparam \in_data_shunt~7 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][5] (
	.clk(clk),
	.d(\in_data_shunt~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][5]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][5] .is_wysiwyg = "true";
defparam \in_data_shunt[0][5] .power_up = "low";

cycloneiv_lcell_comb \source_data~7 (
	.dataa(in_data[5]),
	.datab(\in_data_shunt[0][5]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~7_combout ),
	.cout());
defparam \source_data~7 .lut_mask = 16'hAACC;
defparam \source_data~7 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][6] (
	.clk(clk),
	.d(in_data[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][6]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][6] .is_wysiwyg = "true";
defparam \in_data_shunt[1][6] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~8 (
	.dataa(in_data[6]),
	.datab(\in_data_shunt[1][6]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~8_combout ),
	.cout());
defparam \in_data_shunt~8 .lut_mask = 16'hAACC;
defparam \in_data_shunt~8 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][6] (
	.clk(clk),
	.d(\in_data_shunt~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][6]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][6] .is_wysiwyg = "true";
defparam \in_data_shunt[0][6] .power_up = "low";

cycloneiv_lcell_comb \source_data~8 (
	.dataa(in_data[6]),
	.datab(\in_data_shunt[0][6]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~8_combout ),
	.cout());
defparam \source_data~8 .lut_mask = 16'hAACC;
defparam \source_data~8 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][7] (
	.clk(clk),
	.d(in_data[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][7]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][7] .is_wysiwyg = "true";
defparam \in_data_shunt[1][7] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~9 (
	.dataa(in_data[7]),
	.datab(\in_data_shunt[1][7]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~9_combout ),
	.cout());
defparam \in_data_shunt~9 .lut_mask = 16'hAACC;
defparam \in_data_shunt~9 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][7] (
	.clk(clk),
	.d(\in_data_shunt~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][7]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][7] .is_wysiwyg = "true";
defparam \in_data_shunt[0][7] .power_up = "low";

cycloneiv_lcell_comb \source_data~9 (
	.dataa(in_data[7]),
	.datab(\in_data_shunt[0][7]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~9_combout ),
	.cout());
defparam \source_data~9 .lut_mask = 16'hAACC;
defparam \source_data~9 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][8] (
	.clk(clk),
	.d(in_data[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][8]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][8] .is_wysiwyg = "true";
defparam \in_data_shunt[1][8] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~10 (
	.dataa(in_data[8]),
	.datab(\in_data_shunt[1][8]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~10_combout ),
	.cout());
defparam \in_data_shunt~10 .lut_mask = 16'hAACC;
defparam \in_data_shunt~10 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][8] (
	.clk(clk),
	.d(\in_data_shunt~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][8]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][8] .is_wysiwyg = "true";
defparam \in_data_shunt[0][8] .power_up = "low";

cycloneiv_lcell_comb \source_data~10 (
	.dataa(in_data[8]),
	.datab(\in_data_shunt[0][8]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~10_combout ),
	.cout());
defparam \source_data~10 .lut_mask = 16'hAACC;
defparam \source_data~10 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][9] (
	.clk(clk),
	.d(in_data[9]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][9]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][9] .is_wysiwyg = "true";
defparam \in_data_shunt[1][9] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~11 (
	.dataa(in_data[9]),
	.datab(\in_data_shunt[1][9]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~11_combout ),
	.cout());
defparam \in_data_shunt~11 .lut_mask = 16'hAACC;
defparam \in_data_shunt~11 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][9] (
	.clk(clk),
	.d(\in_data_shunt~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][9]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][9] .is_wysiwyg = "true";
defparam \in_data_shunt[0][9] .power_up = "low";

cycloneiv_lcell_comb \source_data~11 (
	.dataa(in_data[9]),
	.datab(\in_data_shunt[0][9]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~11_combout ),
	.cout());
defparam \source_data~11 .lut_mask = 16'hAACC;
defparam \source_data~11 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][10] (
	.clk(clk),
	.d(in_data[10]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][10]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][10] .is_wysiwyg = "true";
defparam \in_data_shunt[1][10] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~12 (
	.dataa(in_data[10]),
	.datab(\in_data_shunt[1][10]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~12_combout ),
	.cout());
defparam \in_data_shunt~12 .lut_mask = 16'hAACC;
defparam \in_data_shunt~12 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][10] (
	.clk(clk),
	.d(\in_data_shunt~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][10]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][10] .is_wysiwyg = "true";
defparam \in_data_shunt[0][10] .power_up = "low";

cycloneiv_lcell_comb \source_data~12 (
	.dataa(in_data[10]),
	.datab(\in_data_shunt[0][10]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~12_combout ),
	.cout());
defparam \source_data~12 .lut_mask = 16'hAACC;
defparam \source_data~12 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][11] (
	.clk(clk),
	.d(in_data[11]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][11]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][11] .is_wysiwyg = "true";
defparam \in_data_shunt[1][11] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~13 (
	.dataa(in_data[11]),
	.datab(\in_data_shunt[1][11]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~13_combout ),
	.cout());
defparam \in_data_shunt~13 .lut_mask = 16'hAACC;
defparam \in_data_shunt~13 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][11] (
	.clk(clk),
	.d(\in_data_shunt~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][11]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][11] .is_wysiwyg = "true";
defparam \in_data_shunt[0][11] .power_up = "low";

cycloneiv_lcell_comb \source_data~13 (
	.dataa(in_data[11]),
	.datab(\in_data_shunt[0][11]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~13_combout ),
	.cout());
defparam \source_data~13 .lut_mask = 16'hAACC;
defparam \source_data~13 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][12] (
	.clk(clk),
	.d(in_data[12]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][12]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][12] .is_wysiwyg = "true";
defparam \in_data_shunt[1][12] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~14 (
	.dataa(in_data[12]),
	.datab(\in_data_shunt[1][12]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~14_combout ),
	.cout());
defparam \in_data_shunt~14 .lut_mask = 16'hAACC;
defparam \in_data_shunt~14 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][12] (
	.clk(clk),
	.d(\in_data_shunt~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][12]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][12] .is_wysiwyg = "true";
defparam \in_data_shunt[0][12] .power_up = "low";

cycloneiv_lcell_comb \source_data~14 (
	.dataa(in_data[12]),
	.datab(\in_data_shunt[0][12]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~14_combout ),
	.cout());
defparam \source_data~14 .lut_mask = 16'hAACC;
defparam \source_data~14 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][13] (
	.clk(clk),
	.d(in_data[13]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][13]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][13] .is_wysiwyg = "true";
defparam \in_data_shunt[1][13] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~15 (
	.dataa(in_data[13]),
	.datab(\in_data_shunt[1][13]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~15_combout ),
	.cout());
defparam \in_data_shunt~15 .lut_mask = 16'hAACC;
defparam \in_data_shunt~15 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][13] (
	.clk(clk),
	.d(\in_data_shunt~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][13]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][13] .is_wysiwyg = "true";
defparam \in_data_shunt[0][13] .power_up = "low";

cycloneiv_lcell_comb \source_data~15 (
	.dataa(in_data[13]),
	.datab(\in_data_shunt[0][13]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~15_combout ),
	.cout());
defparam \source_data~15 .lut_mask = 16'hAACC;
defparam \source_data~15 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][14] (
	.clk(clk),
	.d(in_data[14]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][14]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][14] .is_wysiwyg = "true";
defparam \in_data_shunt[1][14] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~16 (
	.dataa(in_data[14]),
	.datab(\in_data_shunt[1][14]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~16_combout ),
	.cout());
defparam \in_data_shunt~16 .lut_mask = 16'hAACC;
defparam \in_data_shunt~16 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][14] (
	.clk(clk),
	.d(\in_data_shunt~16_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][14]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][14] .is_wysiwyg = "true";
defparam \in_data_shunt[0][14] .power_up = "low";

cycloneiv_lcell_comb \source_data~16 (
	.dataa(in_data[14]),
	.datab(\in_data_shunt[0][14]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~16_combout ),
	.cout());
defparam \source_data~16 .lut_mask = 16'hAACC;
defparam \source_data~16 .sum_lutc_input = "datac";

dffeas \in_data_shunt[1][15] (
	.clk(clk),
	.d(in_data[15]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\shunt_p~2_combout ),
	.q(\in_data_shunt[1][15]~q ),
	.prn(vcc));
defparam \in_data_shunt[1][15] .is_wysiwyg = "true";
defparam \in_data_shunt[1][15] .power_up = "low";

cycloneiv_lcell_comb \in_data_shunt~17 (
	.dataa(in_data[15]),
	.datab(\in_data_shunt[1][15]~q ),
	.datac(gnd),
	.datad(\shunt_p~1_combout ),
	.cin(gnd),
	.combout(\in_data_shunt~17_combout ),
	.cout());
defparam \in_data_shunt~17 .lut_mask = 16'hAACC;
defparam \in_data_shunt~17 .sum_lutc_input = "datac";

dffeas \in_data_shunt[0][15] (
	.clk(clk),
	.d(\in_data_shunt~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_data_shunt[0][4]~2_combout ),
	.q(\in_data_shunt[0][15]~q ),
	.prn(vcc));
defparam \in_data_shunt[0][15] .is_wysiwyg = "true";
defparam \in_data_shunt[0][15] .power_up = "low";

cycloneiv_lcell_comb \source_data~17 (
	.dataa(in_data[15]),
	.datab(\in_data_shunt[0][15]~q ),
	.datac(gnd),
	.datad(\out_data_p~1_combout ),
	.cin(gnd),
	.combout(\source_data~17_combout ),
	.cout());
defparam \source_data~17 .lut_mask = 16'hAACC;
defparam \source_data~17 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_bit_reverse_core (
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	out_stall,
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Add0,
	Add01,
	rd_valid_dd1,
	out_stall_d1,
	rd_enable,
	out_valid,
	out_enable,
	rd_valid1,
	processing_while_write1,
	out_valid1,
	out_real_0,
	out_real_1,
	out_real_2,
	out_real_3,
	out_real_4,
	out_real_5,
	out_real_6,
	out_real_7,
	out_imag_0,
	out_imag_1,
	out_imag_2,
	out_imag_3,
	out_imag_4,
	out_imag_5,
	out_imag_6,
	out_imag_7,
	out_valid2,
	out_valid3,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	out_stall;
input 	curr_blk_s_2;
input 	curr_blk_s_1;
input 	curr_blk_s_0;
input 	curr_blk_s_3;
input 	Add0;
input 	Add01;
output 	rd_valid_dd1;
output 	out_stall_d1;
output 	rd_enable;
input 	out_valid;
input 	out_enable;
output 	rd_valid1;
output 	processing_while_write1;
input 	out_valid1;
input 	out_real_0;
input 	out_real_1;
input 	out_real_2;
input 	out_real_3;
input 	out_real_4;
input 	out_real_5;
input 	out_real_6;
input 	out_real_7;
input 	out_imag_0;
input 	out_imag_1;
input 	out_imag_2;
input 	out_imag_3;
input 	out_imag_4;
input 	out_imag_5;
input 	out_imag_6;
input 	out_imag_7;
output 	out_valid2;
output 	out_valid3;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \wr_addr_inst|addr_s[0]~q ;
wire \wr_addr_inst|addr_s[2]~q ;
wire \wr_addr_inst|addr_s[1]~q ;
wire \wr_addr_inst|Equal0~1_combout ;
wire \rd_addr_inst|addr_s[0]~q ;
wire \rd_addr_inst|addr_s[1]~q ;
wire \rd_addr_inst|addr_s[2]~q ;
wire \rd_addr_inst|Equal0~1_combout ;
wire \indexing~q ;
wire \indexing~0_combout ;
wire \between_datasets_p~0_combout ;
wire \between_datasets~q ;
wire \rd_enable~1_combout ;
wire \rd_enable~2_combout ;
wire \rd_valid_d~q ;
wire \rd_valid~0_combout ;
wire \rd_valid~1_combout ;


ifft_8p_auk_dspip_bit_reverse_addr_control rd_addr_inst(
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Add0(Add0),
	.Add01(Add01),
	.rd_valid(rd_valid1),
	.rd_enable(\rd_enable~2_combout ),
	.addr_s_0(\rd_addr_inst|addr_s[0]~q ),
	.addr_s_1(\rd_addr_inst|addr_s[1]~q ),
	.addr_s_2(\rd_addr_inst|addr_s[2]~q ),
	.Equal0(\rd_addr_inst|Equal0~1_combout ),
	.indexing(\indexing~q ),
	.clk(clk),
	.reset(reset));

ifft_8p_altera_fft_dual_port_ram real_buf(
	.q_b_8(q_b_8),
	.q_b_9(q_b_9),
	.q_b_10(q_b_10),
	.q_b_11(q_b_11),
	.q_b_12(q_b_12),
	.q_b_13(q_b_13),
	.q_b_14(q_b_14),
	.q_b_15(q_b_15),
	.q_b_0(q_b_0),
	.q_b_1(q_b_1),
	.q_b_2(q_b_2),
	.q_b_3(q_b_3),
	.q_b_4(q_b_4),
	.q_b_5(q_b_5),
	.q_b_6(q_b_6),
	.q_b_7(q_b_7),
	.out_valid(out_valid1),
	.addr_s_0(\wr_addr_inst|addr_s[0]~q ),
	.addr_s_2(\wr_addr_inst|addr_s[2]~q ),
	.addr_s_1(\wr_addr_inst|addr_s[1]~q ),
	.out_real_0(out_real_0),
	.addr_s_01(\rd_addr_inst|addr_s[0]~q ),
	.addr_s_11(\rd_addr_inst|addr_s[1]~q ),
	.addr_s_21(\rd_addr_inst|addr_s[2]~q ),
	.out_real_1(out_real_1),
	.out_real_2(out_real_2),
	.out_real_3(out_real_3),
	.out_real_4(out_real_4),
	.out_real_5(out_real_5),
	.out_real_6(out_real_6),
	.out_real_7(out_real_7),
	.out_imag_0(out_imag_0),
	.out_imag_1(out_imag_1),
	.out_imag_2(out_imag_2),
	.out_imag_3(out_imag_3),
	.out_imag_4(out_imag_4),
	.out_imag_5(out_imag_5),
	.out_imag_6(out_imag_6),
	.out_imag_7(out_imag_7),
	.out_valid1(out_valid2),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_bit_reverse_addr_control_1 wr_addr_inst(
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_1(curr_blk_s_1),
	.curr_blk_s_0(curr_blk_s_0),
	.curr_blk_s_3(curr_blk_s_3),
	.Add0(Add0),
	.Add01(Add01),
	.out_valid(out_valid1),
	.addr_s_0(\wr_addr_inst|addr_s[0]~q ),
	.addr_s_2(\wr_addr_inst|addr_s[2]~q ),
	.addr_s_1(\wr_addr_inst|addr_s[1]~q ),
	.Equal0(\wr_addr_inst|Equal0~1_combout ),
	.indexing(\indexing~q ),
	.clk(clk),
	.reset(reset));

dffeas indexing(
	.clk(clk),
	.d(\indexing~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\indexing~q ),
	.prn(vcc));
defparam indexing.is_wysiwyg = "true";
defparam indexing.power_up = "low";

cycloneiv_lcell_comb \indexing~0 (
	.dataa(gnd),
	.datab(\indexing~q ),
	.datac(out_valid1),
	.datad(\wr_addr_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\indexing~0_combout ),
	.cout());
defparam \indexing~0 .lut_mask = 16'hC33C;
defparam \indexing~0 .sum_lutc_input = "datac";

dffeas rd_valid_dd(
	.clk(clk),
	.d(\rd_valid_d~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_enable~2_combout ),
	.q(rd_valid_dd1),
	.prn(vcc));
defparam rd_valid_dd.is_wysiwyg = "true";
defparam rd_valid_dd.power_up = "low";

dffeas out_stall_d(
	.clk(clk),
	.d(out_stall),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_stall_d1),
	.prn(vcc));
defparam out_stall_d.is_wysiwyg = "true";
defparam out_stall_d.power_up = "low";

cycloneiv_lcell_comb \rd_enable~0 (
	.dataa(\between_datasets~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(out_stall_d1),
	.cin(gnd),
	.combout(rd_enable),
	.cout());
defparam \rd_enable~0 .lut_mask = 16'hAAFF;
defparam \rd_enable~0 .sum_lutc_input = "datac";

dffeas rd_valid(
	.clk(clk),
	.d(\rd_valid~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(rd_valid1),
	.prn(vcc));
defparam rd_valid.is_wysiwyg = "true";
defparam rd_valid.power_up = "low";

dffeas processing_while_write(
	.clk(clk),
	.d(\wr_addr_inst|Equal0~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid1),
	.q(processing_while_write1),
	.prn(vcc));
defparam processing_while_write.is_wysiwyg = "true";
defparam processing_while_write.power_up = "low";

cycloneiv_lcell_comb \out_valid~4 (
	.dataa(\between_datasets~q ),
	.datab(out_stall_d1),
	.datac(out_valid),
	.datad(out_enable),
	.cin(gnd),
	.combout(out_valid2),
	.cout());
defparam \out_valid~4 .lut_mask = 16'hFFFB;
defparam \out_valid~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_valid~5 (
	.dataa(\between_datasets~q ),
	.datab(out_stall_d1),
	.datac(rd_valid_dd1),
	.datad(out_valid1),
	.cin(gnd),
	.combout(out_valid3),
	.cout());
defparam \out_valid~5 .lut_mask = 16'hFFFB;
defparam \out_valid~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \between_datasets_p~0 (
	.dataa(out_valid1),
	.datab(\wr_addr_inst|Equal0~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\between_datasets_p~0_combout ),
	.cout());
defparam \between_datasets_p~0 .lut_mask = 16'hBBBB;
defparam \between_datasets_p~0 .sum_lutc_input = "datac";

dffeas between_datasets(
	.clk(clk),
	.d(\between_datasets_p~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid1),
	.q(\between_datasets~q ),
	.prn(vcc));
defparam between_datasets.is_wysiwyg = "true";
defparam between_datasets.power_up = "low";

cycloneiv_lcell_comb \rd_enable~1 (
	.dataa(\wr_addr_inst|addr_s[0]~q ),
	.datab(\wr_addr_inst|addr_s[2]~q ),
	.datac(\wr_addr_inst|addr_s[1]~q ),
	.datad(\between_datasets~q ),
	.cin(gnd),
	.combout(\rd_enable~1_combout ),
	.cout());
defparam \rd_enable~1 .lut_mask = 16'h7FFF;
defparam \rd_enable~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \rd_enable~2 (
	.dataa(rd_enable),
	.datab(out_valid),
	.datac(\rd_enable~1_combout ),
	.datad(out_enable),
	.cin(gnd),
	.combout(\rd_enable~2_combout ),
	.cout());
defparam \rd_enable~2 .lut_mask = 16'hFFFE;
defparam \rd_enable~2 .sum_lutc_input = "datac";

dffeas rd_valid_d(
	.clk(clk),
	.d(rd_valid1),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\rd_enable~2_combout ),
	.q(\rd_valid_d~q ),
	.prn(vcc));
defparam rd_valid_d.is_wysiwyg = "true";
defparam rd_valid_d.power_up = "low";

cycloneiv_lcell_comb \rd_valid~0 (
	.dataa(rd_valid1),
	.datab(out_valid1),
	.datac(\wr_addr_inst|Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\rd_valid~0_combout ),
	.cout());
defparam \rd_valid~0 .lut_mask = 16'hEFEF;
defparam \rd_valid~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \rd_valid~1 (
	.dataa(\rd_valid~0_combout ),
	.datab(\wr_addr_inst|Equal0~1_combout ),
	.datac(\rd_enable~2_combout ),
	.datad(\rd_addr_inst|Equal0~1_combout ),
	.cin(gnd),
	.combout(\rd_valid~1_combout ),
	.cout());
defparam \rd_valid~1 .lut_mask = 16'hBFFF;
defparam \rd_valid~1 .sum_lutc_input = "datac";

endmodule

module ifft_8p_altera_fft_dual_port_ram (
	q_b_8,
	q_b_9,
	q_b_10,
	q_b_11,
	q_b_12,
	q_b_13,
	q_b_14,
	q_b_15,
	q_b_0,
	q_b_1,
	q_b_2,
	q_b_3,
	q_b_4,
	q_b_5,
	q_b_6,
	q_b_7,
	out_valid,
	addr_s_0,
	addr_s_2,
	addr_s_1,
	out_real_0,
	addr_s_01,
	addr_s_11,
	addr_s_21,
	out_real_1,
	out_real_2,
	out_real_3,
	out_real_4,
	out_real_5,
	out_real_6,
	out_real_7,
	out_imag_0,
	out_imag_1,
	out_imag_2,
	out_imag_3,
	out_imag_4,
	out_imag_5,
	out_imag_6,
	out_imag_7,
	out_valid1,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	q_b_8;
output 	q_b_9;
output 	q_b_10;
output 	q_b_11;
output 	q_b_12;
output 	q_b_13;
output 	q_b_14;
output 	q_b_15;
output 	q_b_0;
output 	q_b_1;
output 	q_b_2;
output 	q_b_3;
output 	q_b_4;
output 	q_b_5;
output 	q_b_6;
output 	q_b_7;
input 	out_valid;
input 	addr_s_0;
input 	addr_s_2;
input 	addr_s_1;
input 	out_real_0;
input 	addr_s_01;
input 	addr_s_11;
input 	addr_s_21;
input 	out_real_1;
input 	out_real_2;
input 	out_real_3;
input 	out_real_4;
input 	out_real_5;
input 	out_real_6;
input 	out_real_7;
input 	out_imag_0;
input 	out_imag_1;
input 	out_imag_2;
input 	out_imag_3;
input 	out_imag_4;
input 	out_imag_5;
input 	out_imag_6;
input 	out_imag_7;
input 	out_valid1;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altsyncram_1 \old_ram_gen:old_ram_component (
	.q_b({q_b_15,q_b_14,q_b_13,q_b_12,q_b_11,q_b_10,q_b_9,q_b_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.wren_a(out_valid),
	.address_a({addr_s_2,addr_s_1,addr_s_0}),
	.data_a({out_real_7,out_real_6,out_real_5,out_real_4,out_real_3,out_real_2,out_real_1,out_real_0,out_imag_7,out_imag_6,out_imag_5,out_imag_4,out_imag_3,out_imag_2,out_imag_1,out_imag_0}),
	.address_b({addr_s_21,addr_s_11,addr_s_01}),
	.clocken0(out_valid1),
	.clock0(clk),
	.aclr0(reset_n));

endmodule

module ifft_8p_altsyncram_1 (
	q_b,
	wren_a,
	address_a,
	data_a,
	address_b,
	clocken0,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[2:0] address_a;
input 	[15:0] data_a;
input 	[2:0] address_b;
input 	clocken0;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altsyncram_k9p3 auto_generated(
	.q_b({q_b[15],q_b[14],q_b[13],q_b[12],q_b[11],q_b[10],q_b[9],q_b[8],q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.wren_a(wren_a),
	.address_a({address_a[2],address_a[1],address_a[0]}),
	.data_a({data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_b({address_b[2],address_b[1],address_b[0]}),
	.clocken0(clocken0),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_altsyncram_k9p3 (
	q_b,
	wren_a,
	address_a,
	data_a,
	address_b,
	clocken0,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_b;
input 	wren_a;
input 	[2:0] address_a;
input 	[15:0] data_a;
input 	[2:0] address_b;
input 	clocken0;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a8_PORTBDATAOUT_bus;
wire [143:0] ram_block1a9_PORTBDATAOUT_bus;
wire [143:0] ram_block1a10_PORTBDATAOUT_bus;
wire [143:0] ram_block1a11_PORTBDATAOUT_bus;
wire [143:0] ram_block1a12_PORTBDATAOUT_bus;
wire [143:0] ram_block1a13_PORTBDATAOUT_bus;
wire [143:0] ram_block1a14_PORTBDATAOUT_bus;
wire [143:0] ram_block1a15_PORTBDATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_b[8] = ram_block1a8_PORTBDATAOUT_bus[0];

assign q_b[9] = ram_block1a9_PORTBDATAOUT_bus[0];

assign q_b[10] = ram_block1a10_PORTBDATAOUT_bus[0];

assign q_b[11] = ram_block1a11_PORTBDATAOUT_bus[0];

assign q_b[12] = ram_block1a12_PORTBDATAOUT_bus[0];

assign q_b[13] = ram_block1a13_PORTBDATAOUT_bus[0];

assign q_b[14] = ram_block1a14_PORTBDATAOUT_bus[0];

assign q_b[15] = ram_block1a15_PORTBDATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneiv_ram_block ram_block1a8(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[8]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a8_PORTBDATAOUT_bus));
defparam ram_block1a8.clk0_core_clock_enable = "ena0";
defparam ram_block1a8.clk0_input_clock_enable = "ena0";
defparam ram_block1a8.clk0_output_clock_enable = "ena0";
defparam ram_block1a8.data_interleave_offset_in_bits = 1;
defparam ram_block1a8.data_interleave_width_in_bits = 1;
defparam ram_block1a8.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a8.mixed_port_feed_through_mode = "old";
defparam ram_block1a8.operation_mode = "dual_port";
defparam ram_block1a8.port_a_address_clear = "none";
defparam ram_block1a8.port_a_address_width = 3;
defparam ram_block1a8.port_a_data_out_clear = "none";
defparam ram_block1a8.port_a_data_out_clock = "none";
defparam ram_block1a8.port_a_data_width = 1;
defparam ram_block1a8.port_a_first_address = 0;
defparam ram_block1a8.port_a_first_bit_number = 8;
defparam ram_block1a8.port_a_last_address = 7;
defparam ram_block1a8.port_a_logical_ram_depth = 8;
defparam ram_block1a8.port_a_logical_ram_width = 16;
defparam ram_block1a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_address_clear = "clear0";
defparam ram_block1a8.port_b_address_clock = "clock0";
defparam ram_block1a8.port_b_address_width = 3;
defparam ram_block1a8.port_b_data_out_clear = "clear0";
defparam ram_block1a8.port_b_data_out_clock = "clock0";
defparam ram_block1a8.port_b_data_width = 1;
defparam ram_block1a8.port_b_first_address = 0;
defparam ram_block1a8.port_b_first_bit_number = 8;
defparam ram_block1a8.port_b_last_address = 7;
defparam ram_block1a8.port_b_logical_ram_depth = 8;
defparam ram_block1a8.port_b_logical_ram_width = 16;
defparam ram_block1a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a8.port_b_read_enable_clock = "clock0";
defparam ram_block1a8.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a9(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[9]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a9_PORTBDATAOUT_bus));
defparam ram_block1a9.clk0_core_clock_enable = "ena0";
defparam ram_block1a9.clk0_input_clock_enable = "ena0";
defparam ram_block1a9.clk0_output_clock_enable = "ena0";
defparam ram_block1a9.data_interleave_offset_in_bits = 1;
defparam ram_block1a9.data_interleave_width_in_bits = 1;
defparam ram_block1a9.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a9.mixed_port_feed_through_mode = "old";
defparam ram_block1a9.operation_mode = "dual_port";
defparam ram_block1a9.port_a_address_clear = "none";
defparam ram_block1a9.port_a_address_width = 3;
defparam ram_block1a9.port_a_data_out_clear = "none";
defparam ram_block1a9.port_a_data_out_clock = "none";
defparam ram_block1a9.port_a_data_width = 1;
defparam ram_block1a9.port_a_first_address = 0;
defparam ram_block1a9.port_a_first_bit_number = 9;
defparam ram_block1a9.port_a_last_address = 7;
defparam ram_block1a9.port_a_logical_ram_depth = 8;
defparam ram_block1a9.port_a_logical_ram_width = 16;
defparam ram_block1a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_address_clear = "clear0";
defparam ram_block1a9.port_b_address_clock = "clock0";
defparam ram_block1a9.port_b_address_width = 3;
defparam ram_block1a9.port_b_data_out_clear = "clear0";
defparam ram_block1a9.port_b_data_out_clock = "clock0";
defparam ram_block1a9.port_b_data_width = 1;
defparam ram_block1a9.port_b_first_address = 0;
defparam ram_block1a9.port_b_first_bit_number = 9;
defparam ram_block1a9.port_b_last_address = 7;
defparam ram_block1a9.port_b_logical_ram_depth = 8;
defparam ram_block1a9.port_b_logical_ram_width = 16;
defparam ram_block1a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a9.port_b_read_enable_clock = "clock0";
defparam ram_block1a9.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a10(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[10]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a10_PORTBDATAOUT_bus));
defparam ram_block1a10.clk0_core_clock_enable = "ena0";
defparam ram_block1a10.clk0_input_clock_enable = "ena0";
defparam ram_block1a10.clk0_output_clock_enable = "ena0";
defparam ram_block1a10.data_interleave_offset_in_bits = 1;
defparam ram_block1a10.data_interleave_width_in_bits = 1;
defparam ram_block1a10.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a10.mixed_port_feed_through_mode = "old";
defparam ram_block1a10.operation_mode = "dual_port";
defparam ram_block1a10.port_a_address_clear = "none";
defparam ram_block1a10.port_a_address_width = 3;
defparam ram_block1a10.port_a_data_out_clear = "none";
defparam ram_block1a10.port_a_data_out_clock = "none";
defparam ram_block1a10.port_a_data_width = 1;
defparam ram_block1a10.port_a_first_address = 0;
defparam ram_block1a10.port_a_first_bit_number = 10;
defparam ram_block1a10.port_a_last_address = 7;
defparam ram_block1a10.port_a_logical_ram_depth = 8;
defparam ram_block1a10.port_a_logical_ram_width = 16;
defparam ram_block1a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_address_clear = "clear0";
defparam ram_block1a10.port_b_address_clock = "clock0";
defparam ram_block1a10.port_b_address_width = 3;
defparam ram_block1a10.port_b_data_out_clear = "clear0";
defparam ram_block1a10.port_b_data_out_clock = "clock0";
defparam ram_block1a10.port_b_data_width = 1;
defparam ram_block1a10.port_b_first_address = 0;
defparam ram_block1a10.port_b_first_bit_number = 10;
defparam ram_block1a10.port_b_last_address = 7;
defparam ram_block1a10.port_b_logical_ram_depth = 8;
defparam ram_block1a10.port_b_logical_ram_width = 16;
defparam ram_block1a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a10.port_b_read_enable_clock = "clock0";
defparam ram_block1a10.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a11(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[11]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a11_PORTBDATAOUT_bus));
defparam ram_block1a11.clk0_core_clock_enable = "ena0";
defparam ram_block1a11.clk0_input_clock_enable = "ena0";
defparam ram_block1a11.clk0_output_clock_enable = "ena0";
defparam ram_block1a11.data_interleave_offset_in_bits = 1;
defparam ram_block1a11.data_interleave_width_in_bits = 1;
defparam ram_block1a11.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a11.mixed_port_feed_through_mode = "old";
defparam ram_block1a11.operation_mode = "dual_port";
defparam ram_block1a11.port_a_address_clear = "none";
defparam ram_block1a11.port_a_address_width = 3;
defparam ram_block1a11.port_a_data_out_clear = "none";
defparam ram_block1a11.port_a_data_out_clock = "none";
defparam ram_block1a11.port_a_data_width = 1;
defparam ram_block1a11.port_a_first_address = 0;
defparam ram_block1a11.port_a_first_bit_number = 11;
defparam ram_block1a11.port_a_last_address = 7;
defparam ram_block1a11.port_a_logical_ram_depth = 8;
defparam ram_block1a11.port_a_logical_ram_width = 16;
defparam ram_block1a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_address_clear = "clear0";
defparam ram_block1a11.port_b_address_clock = "clock0";
defparam ram_block1a11.port_b_address_width = 3;
defparam ram_block1a11.port_b_data_out_clear = "clear0";
defparam ram_block1a11.port_b_data_out_clock = "clock0";
defparam ram_block1a11.port_b_data_width = 1;
defparam ram_block1a11.port_b_first_address = 0;
defparam ram_block1a11.port_b_first_bit_number = 11;
defparam ram_block1a11.port_b_last_address = 7;
defparam ram_block1a11.port_b_logical_ram_depth = 8;
defparam ram_block1a11.port_b_logical_ram_width = 16;
defparam ram_block1a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a11.port_b_read_enable_clock = "clock0";
defparam ram_block1a11.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a12(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[12]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a12_PORTBDATAOUT_bus));
defparam ram_block1a12.clk0_core_clock_enable = "ena0";
defparam ram_block1a12.clk0_input_clock_enable = "ena0";
defparam ram_block1a12.clk0_output_clock_enable = "ena0";
defparam ram_block1a12.data_interleave_offset_in_bits = 1;
defparam ram_block1a12.data_interleave_width_in_bits = 1;
defparam ram_block1a12.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a12.mixed_port_feed_through_mode = "old";
defparam ram_block1a12.operation_mode = "dual_port";
defparam ram_block1a12.port_a_address_clear = "none";
defparam ram_block1a12.port_a_address_width = 3;
defparam ram_block1a12.port_a_data_out_clear = "none";
defparam ram_block1a12.port_a_data_out_clock = "none";
defparam ram_block1a12.port_a_data_width = 1;
defparam ram_block1a12.port_a_first_address = 0;
defparam ram_block1a12.port_a_first_bit_number = 12;
defparam ram_block1a12.port_a_last_address = 7;
defparam ram_block1a12.port_a_logical_ram_depth = 8;
defparam ram_block1a12.port_a_logical_ram_width = 16;
defparam ram_block1a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_address_clear = "clear0";
defparam ram_block1a12.port_b_address_clock = "clock0";
defparam ram_block1a12.port_b_address_width = 3;
defparam ram_block1a12.port_b_data_out_clear = "clear0";
defparam ram_block1a12.port_b_data_out_clock = "clock0";
defparam ram_block1a12.port_b_data_width = 1;
defparam ram_block1a12.port_b_first_address = 0;
defparam ram_block1a12.port_b_first_bit_number = 12;
defparam ram_block1a12.port_b_last_address = 7;
defparam ram_block1a12.port_b_logical_ram_depth = 8;
defparam ram_block1a12.port_b_logical_ram_width = 16;
defparam ram_block1a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a12.port_b_read_enable_clock = "clock0";
defparam ram_block1a12.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a13(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[13]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a13_PORTBDATAOUT_bus));
defparam ram_block1a13.clk0_core_clock_enable = "ena0";
defparam ram_block1a13.clk0_input_clock_enable = "ena0";
defparam ram_block1a13.clk0_output_clock_enable = "ena0";
defparam ram_block1a13.data_interleave_offset_in_bits = 1;
defparam ram_block1a13.data_interleave_width_in_bits = 1;
defparam ram_block1a13.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a13.mixed_port_feed_through_mode = "old";
defparam ram_block1a13.operation_mode = "dual_port";
defparam ram_block1a13.port_a_address_clear = "none";
defparam ram_block1a13.port_a_address_width = 3;
defparam ram_block1a13.port_a_data_out_clear = "none";
defparam ram_block1a13.port_a_data_out_clock = "none";
defparam ram_block1a13.port_a_data_width = 1;
defparam ram_block1a13.port_a_first_address = 0;
defparam ram_block1a13.port_a_first_bit_number = 13;
defparam ram_block1a13.port_a_last_address = 7;
defparam ram_block1a13.port_a_logical_ram_depth = 8;
defparam ram_block1a13.port_a_logical_ram_width = 16;
defparam ram_block1a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_address_clear = "clear0";
defparam ram_block1a13.port_b_address_clock = "clock0";
defparam ram_block1a13.port_b_address_width = 3;
defparam ram_block1a13.port_b_data_out_clear = "clear0";
defparam ram_block1a13.port_b_data_out_clock = "clock0";
defparam ram_block1a13.port_b_data_width = 1;
defparam ram_block1a13.port_b_first_address = 0;
defparam ram_block1a13.port_b_first_bit_number = 13;
defparam ram_block1a13.port_b_last_address = 7;
defparam ram_block1a13.port_b_logical_ram_depth = 8;
defparam ram_block1a13.port_b_logical_ram_width = 16;
defparam ram_block1a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a13.port_b_read_enable_clock = "clock0";
defparam ram_block1a13.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a14(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[14]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a14_PORTBDATAOUT_bus));
defparam ram_block1a14.clk0_core_clock_enable = "ena0";
defparam ram_block1a14.clk0_input_clock_enable = "ena0";
defparam ram_block1a14.clk0_output_clock_enable = "ena0";
defparam ram_block1a14.data_interleave_offset_in_bits = 1;
defparam ram_block1a14.data_interleave_width_in_bits = 1;
defparam ram_block1a14.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a14.mixed_port_feed_through_mode = "old";
defparam ram_block1a14.operation_mode = "dual_port";
defparam ram_block1a14.port_a_address_clear = "none";
defparam ram_block1a14.port_a_address_width = 3;
defparam ram_block1a14.port_a_data_out_clear = "none";
defparam ram_block1a14.port_a_data_out_clock = "none";
defparam ram_block1a14.port_a_data_width = 1;
defparam ram_block1a14.port_a_first_address = 0;
defparam ram_block1a14.port_a_first_bit_number = 14;
defparam ram_block1a14.port_a_last_address = 7;
defparam ram_block1a14.port_a_logical_ram_depth = 8;
defparam ram_block1a14.port_a_logical_ram_width = 16;
defparam ram_block1a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_address_clear = "clear0";
defparam ram_block1a14.port_b_address_clock = "clock0";
defparam ram_block1a14.port_b_address_width = 3;
defparam ram_block1a14.port_b_data_out_clear = "clear0";
defparam ram_block1a14.port_b_data_out_clock = "clock0";
defparam ram_block1a14.port_b_data_width = 1;
defparam ram_block1a14.port_b_first_address = 0;
defparam ram_block1a14.port_b_first_bit_number = 14;
defparam ram_block1a14.port_b_last_address = 7;
defparam ram_block1a14.port_b_logical_ram_depth = 8;
defparam ram_block1a14.port_b_logical_ram_width = 16;
defparam ram_block1a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a14.port_b_read_enable_clock = "clock0";
defparam ram_block1a14.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a15(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[15]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a15_PORTBDATAOUT_bus));
defparam ram_block1a15.clk0_core_clock_enable = "ena0";
defparam ram_block1a15.clk0_input_clock_enable = "ena0";
defparam ram_block1a15.clk0_output_clock_enable = "ena0";
defparam ram_block1a15.data_interleave_offset_in_bits = 1;
defparam ram_block1a15.data_interleave_width_in_bits = 1;
defparam ram_block1a15.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a15.mixed_port_feed_through_mode = "old";
defparam ram_block1a15.operation_mode = "dual_port";
defparam ram_block1a15.port_a_address_clear = "none";
defparam ram_block1a15.port_a_address_width = 3;
defparam ram_block1a15.port_a_data_out_clear = "none";
defparam ram_block1a15.port_a_data_out_clock = "none";
defparam ram_block1a15.port_a_data_width = 1;
defparam ram_block1a15.port_a_first_address = 0;
defparam ram_block1a15.port_a_first_bit_number = 15;
defparam ram_block1a15.port_a_last_address = 7;
defparam ram_block1a15.port_a_logical_ram_depth = 8;
defparam ram_block1a15.port_a_logical_ram_width = 16;
defparam ram_block1a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_address_clear = "clear0";
defparam ram_block1a15.port_b_address_clock = "clock0";
defparam ram_block1a15.port_b_address_width = 3;
defparam ram_block1a15.port_b_data_out_clear = "clear0";
defparam ram_block1a15.port_b_data_out_clock = "clock0";
defparam ram_block1a15.port_b_data_width = 1;
defparam ram_block1a15.port_b_first_address = 0;
defparam ram_block1a15.port_b_first_bit_number = 15;
defparam ram_block1a15.port_b_last_address = 7;
defparam ram_block1a15.port_b_logical_ram_depth = 8;
defparam ram_block1a15.port_b_logical_ram_width = 16;
defparam ram_block1a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a15.port_b_read_enable_clock = "clock0";
defparam ram_block1a15.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a0(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "old";
defparam ram_block1a0.operation_mode = "dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 3;
defparam ram_block1a0.port_a_data_out_clear = "none";
defparam ram_block1a0.port_a_data_out_clock = "none";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 7;
defparam ram_block1a0.port_a_logical_ram_depth = 8;
defparam ram_block1a0.port_a_logical_ram_width = 16;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "clear0";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 3;
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 7;
defparam ram_block1a0.port_b_logical_ram_depth = 8;
defparam ram_block1a0.port_b_logical_ram_width = 16;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a1(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[1]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "old";
defparam ram_block1a1.operation_mode = "dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 3;
defparam ram_block1a1.port_a_data_out_clear = "none";
defparam ram_block1a1.port_a_data_out_clock = "none";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 7;
defparam ram_block1a1.port_a_logical_ram_depth = 8;
defparam ram_block1a1.port_a_logical_ram_width = 16;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "clear0";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 3;
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 7;
defparam ram_block1a1.port_b_logical_ram_depth = 8;
defparam ram_block1a1.port_b_logical_ram_width = 16;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a2(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[2]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "old";
defparam ram_block1a2.operation_mode = "dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 3;
defparam ram_block1a2.port_a_data_out_clear = "none";
defparam ram_block1a2.port_a_data_out_clock = "none";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 7;
defparam ram_block1a2.port_a_logical_ram_depth = 8;
defparam ram_block1a2.port_a_logical_ram_width = 16;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "clear0";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 3;
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 7;
defparam ram_block1a2.port_b_logical_ram_depth = 8;
defparam ram_block1a2.port_b_logical_ram_width = 16;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a3(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[3]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "old";
defparam ram_block1a3.operation_mode = "dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 3;
defparam ram_block1a3.port_a_data_out_clear = "none";
defparam ram_block1a3.port_a_data_out_clock = "none";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 7;
defparam ram_block1a3.port_a_logical_ram_depth = 8;
defparam ram_block1a3.port_a_logical_ram_width = 16;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "clear0";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 3;
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 7;
defparam ram_block1a3.port_b_logical_ram_depth = 8;
defparam ram_block1a3.port_b_logical_ram_width = 16;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a4(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[4]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "old";
defparam ram_block1a4.operation_mode = "dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 3;
defparam ram_block1a4.port_a_data_out_clear = "none";
defparam ram_block1a4.port_a_data_out_clock = "none";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 7;
defparam ram_block1a4.port_a_logical_ram_depth = 8;
defparam ram_block1a4.port_a_logical_ram_width = 16;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "clear0";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 3;
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 7;
defparam ram_block1a4.port_b_logical_ram_depth = 8;
defparam ram_block1a4.port_b_logical_ram_width = 16;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a5(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[5]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "old";
defparam ram_block1a5.operation_mode = "dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 3;
defparam ram_block1a5.port_a_data_out_clear = "none";
defparam ram_block1a5.port_a_data_out_clock = "none";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 7;
defparam ram_block1a5.port_a_logical_ram_depth = 8;
defparam ram_block1a5.port_a_logical_ram_width = 16;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "clear0";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 3;
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 7;
defparam ram_block1a5.port_b_logical_ram_depth = 8;
defparam ram_block1a5.port_b_logical_ram_width = 16;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a6(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[6]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "old";
defparam ram_block1a6.operation_mode = "dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 3;
defparam ram_block1a6.port_a_data_out_clear = "none";
defparam ram_block1a6.port_a_data_out_clock = "none";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 7;
defparam ram_block1a6.port_a_logical_ram_depth = 8;
defparam ram_block1a6.port_a_logical_ram_width = 16;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "clear0";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 3;
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 7;
defparam ram_block1a6.port_b_logical_ram_depth = 8;
defparam ram_block1a6.port_b_logical_ram_width = 16;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";

cycloneiv_ram_block ram_block1a7(
	.portawe(wren_a),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[7]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain(1'b0),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_bit_reverse_core:\\generate_bit_reverse_module:bit_reverse_inst|altera_fft_dual_port_ram:real_buf|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_k9p3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "old";
defparam ram_block1a7.operation_mode = "dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 3;
defparam ram_block1a7.port_a_data_out_clear = "none";
defparam ram_block1a7.port_a_data_out_clock = "none";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 7;
defparam ram_block1a7.port_a_logical_ram_depth = 8;
defparam ram_block1a7.port_a_logical_ram_width = 16;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "clear0";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 3;
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 7;
defparam ram_block1a7.port_b_logical_ram_depth = 8;
defparam ram_block1a7.port_b_logical_ram_width = 16;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";

endmodule

module ifft_8p_auk_dspip_bit_reverse_addr_control (
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Add0,
	Add01,
	rd_valid,
	rd_enable,
	addr_s_0,
	addr_s_1,
	addr_s_2,
	Equal0,
	indexing,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_2;
input 	curr_blk_s_1;
input 	curr_blk_s_0;
input 	curr_blk_s_3;
input 	Add0;
input 	Add01;
input 	rd_valid;
input 	rd_enable;
output 	addr_s_0;
output 	addr_s_1;
output 	addr_s_2;
output 	Equal0;
input 	indexing;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \reverse_carry_adder_inst|cout[1]~0_combout ;
wire \reverse_carry_adder_inst|sum_out[1]~0_combout ;
wire \addr_s~0_combout ;
wire \addr_s~1_combout ;
wire \gen_addr~0_combout ;
wire \Add1~0_combout ;
wire \addr_s~2_combout ;
wire \addr_s~3_combout ;
wire \addr_s~4_combout ;
wire \Equal0~0_combout ;


ifft_8p_auk_dspip_bit_reverse_reverse_carry_adder reverse_carry_adder_inst(
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_3(curr_blk_s_3),
	.addr_s_1(addr_s_1),
	.addr_s_2(addr_s_2),
	.cout_1(\reverse_carry_adder_inst|cout[1]~0_combout ),
	.sum_out_1(\reverse_carry_adder_inst|sum_out[1]~0_combout ));

dffeas \addr_s[0] (
	.clk(clk),
	.d(\addr_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\gen_addr~0_combout ),
	.q(addr_s_0),
	.prn(vcc));
defparam \addr_s[0] .is_wysiwyg = "true";
defparam \addr_s[0] .power_up = "low";

dffeas \addr_s[1] (
	.clk(clk),
	.d(\addr_s~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\gen_addr~0_combout ),
	.q(addr_s_1),
	.prn(vcc));
defparam \addr_s[1] .is_wysiwyg = "true";
defparam \addr_s[1] .power_up = "low";

dffeas \addr_s[2] (
	.clk(clk),
	.d(\addr_s~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\gen_addr~0_combout ),
	.q(addr_s_2),
	.prn(vcc));
defparam \addr_s[2] .is_wysiwyg = "true";
defparam \addr_s[2] .power_up = "low";

cycloneiv_lcell_comb \Equal0~1 (
	.dataa(Add0),
	.datab(\Equal0~0_combout ),
	.datac(Add01),
	.datad(addr_s_2),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hDFFD;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~0 (
	.dataa(indexing),
	.datab(curr_blk_s_1),
	.datac(addr_s_0),
	.datad(\reverse_carry_adder_inst|cout[1]~0_combout ),
	.cin(gnd),
	.combout(\addr_s~0_combout ),
	.cout());
defparam \addr_s~0 .lut_mask = 16'hEBBE;
defparam \addr_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~1 (
	.dataa(\addr_s~0_combout ),
	.datab(indexing),
	.datac(addr_s_0),
	.datad(Equal0),
	.cin(gnd),
	.combout(\addr_s~1_combout ),
	.cout());
defparam \addr_s~1 .lut_mask = 16'hBFFF;
defparam \addr_s~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \gen_addr~0 (
	.dataa(rd_enable),
	.datab(rd_valid),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\gen_addr~0_combout ),
	.cout());
defparam \gen_addr~0 .lut_mask = 16'hEEEE;
defparam \gen_addr~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(addr_s_0),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~2 (
	.dataa(\reverse_carry_adder_inst|sum_out[1]~0_combout ),
	.datab(indexing),
	.datac(\Add1~0_combout ),
	.datad(Equal0),
	.cin(gnd),
	.combout(\addr_s~2_combout ),
	.cout());
defparam \addr_s~2 .lut_mask = 16'hB8FF;
defparam \addr_s~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~3 (
	.dataa(indexing),
	.datab(addr_s_2),
	.datac(addr_s_0),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(\addr_s~3_combout ),
	.cout());
defparam \addr_s~3 .lut_mask = 16'h6996;
defparam \addr_s~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~4 (
	.dataa(curr_blk_s_3),
	.datab(Equal0),
	.datac(indexing),
	.datad(\addr_s~3_combout ),
	.cin(gnd),
	.combout(\addr_s~4_combout ),
	.cout());
defparam \addr_s~4 .lut_mask = 16'hB77B;
defparam \addr_s~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(curr_blk_s_1),
	.datab(addr_s_1),
	.datac(curr_blk_s_0),
	.datad(addr_s_0),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_bit_reverse_reverse_carry_adder (
	curr_blk_s_2,
	curr_blk_s_3,
	addr_s_1,
	addr_s_2,
	cout_1,
	sum_out_1)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_2;
input 	curr_blk_s_3;
input 	addr_s_1;
input 	addr_s_2;
output 	cout_1;
output 	sum_out_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \cout[1]~0 (
	.dataa(addr_s_2),
	.datab(curr_blk_s_3),
	.datac(curr_blk_s_2),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(cout_1),
	.cout());
defparam \cout[1]~0 .lut_mask = 16'hFFFE;
defparam \cout[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \sum_out[1]~0 (
	.dataa(curr_blk_s_3),
	.datab(addr_s_2),
	.datac(curr_blk_s_2),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(sum_out_1),
	.cout());
defparam \sum_out[1]~0 .lut_mask = 16'h6996;
defparam \sum_out[1]~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_bit_reverse_addr_control_1 (
	curr_blk_s_2,
	curr_blk_s_1,
	curr_blk_s_0,
	curr_blk_s_3,
	Add0,
	Add01,
	out_valid,
	addr_s_0,
	addr_s_2,
	addr_s_1,
	Equal0,
	indexing,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_2;
input 	curr_blk_s_1;
input 	curr_blk_s_0;
input 	curr_blk_s_3;
input 	Add0;
input 	Add01;
input 	out_valid;
output 	addr_s_0;
output 	addr_s_2;
output 	addr_s_1;
output 	Equal0;
input 	indexing;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \reverse_carry_adder_inst|cout[1]~0_combout ;
wire \reverse_carry_adder_inst|sum_out[1]~0_combout ;
wire \addr_s~0_combout ;
wire \addr_s~1_combout ;
wire \addr_s~2_combout ;
wire \addr_s~3_combout ;
wire \Add1~0_combout ;
wire \addr_s~4_combout ;
wire \Equal0~0_combout ;


ifft_8p_auk_dspip_bit_reverse_reverse_carry_adder_1 reverse_carry_adder_inst(
	.curr_blk_s_2(curr_blk_s_2),
	.curr_blk_s_3(curr_blk_s_3),
	.addr_s_2(addr_s_2),
	.addr_s_1(addr_s_1),
	.cout_1(\reverse_carry_adder_inst|cout[1]~0_combout ),
	.sum_out_1(\reverse_carry_adder_inst|sum_out[1]~0_combout ));

dffeas \addr_s[0] (
	.clk(clk),
	.d(\addr_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid),
	.q(addr_s_0),
	.prn(vcc));
defparam \addr_s[0] .is_wysiwyg = "true";
defparam \addr_s[0] .power_up = "low";

dffeas \addr_s[2] (
	.clk(clk),
	.d(\addr_s~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid),
	.q(addr_s_2),
	.prn(vcc));
defparam \addr_s[2] .is_wysiwyg = "true";
defparam \addr_s[2] .power_up = "low";

dffeas \addr_s[1] (
	.clk(clk),
	.d(\addr_s~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_valid),
	.q(addr_s_1),
	.prn(vcc));
defparam \addr_s[1] .is_wysiwyg = "true";
defparam \addr_s[1] .power_up = "low";

cycloneiv_lcell_comb \Equal0~1 (
	.dataa(Add0),
	.datab(\Equal0~0_combout ),
	.datac(Add01),
	.datad(addr_s_2),
	.cin(gnd),
	.combout(Equal0),
	.cout());
defparam \Equal0~1 .lut_mask = 16'hBFFB;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~0 (
	.dataa(indexing),
	.datab(curr_blk_s_1),
	.datac(addr_s_0),
	.datad(\reverse_carry_adder_inst|cout[1]~0_combout ),
	.cin(gnd),
	.combout(\addr_s~0_combout ),
	.cout());
defparam \addr_s~0 .lut_mask = 16'hEBBE;
defparam \addr_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~1 (
	.dataa(\addr_s~0_combout ),
	.datab(addr_s_0),
	.datac(Equal0),
	.datad(indexing),
	.cin(gnd),
	.combout(\addr_s~1_combout ),
	.cout());
defparam \addr_s~1 .lut_mask = 16'hFBFF;
defparam \addr_s~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~2 (
	.dataa(indexing),
	.datab(addr_s_2),
	.datac(addr_s_0),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(\addr_s~2_combout ),
	.cout());
defparam \addr_s~2 .lut_mask = 16'h6996;
defparam \addr_s~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~3 (
	.dataa(curr_blk_s_3),
	.datab(Equal0),
	.datac(indexing),
	.datad(\addr_s~2_combout ),
	.cin(gnd),
	.combout(\addr_s~3_combout ),
	.cout());
defparam \addr_s~3 .lut_mask = 16'hEDDE;
defparam \addr_s~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add1~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(addr_s_0),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h0FF0;
defparam \Add1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \addr_s~4 (
	.dataa(\reverse_carry_adder_inst|sum_out[1]~0_combout ),
	.datab(indexing),
	.datac(\Add1~0_combout ),
	.datad(Equal0),
	.cin(gnd),
	.combout(\addr_s~4_combout ),
	.cout());
defparam \addr_s~4 .lut_mask = 16'hFFB8;
defparam \addr_s~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(curr_blk_s_1),
	.datab(addr_s_1),
	.datac(curr_blk_s_0),
	.datad(addr_s_0),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_bit_reverse_reverse_carry_adder_1 (
	curr_blk_s_2,
	curr_blk_s_3,
	addr_s_2,
	addr_s_1,
	cout_1,
	sum_out_1)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_2;
input 	curr_blk_s_3;
input 	addr_s_2;
input 	addr_s_1;
output 	cout_1;
output 	sum_out_1;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



cycloneiv_lcell_comb \cout[1]~0 (
	.dataa(addr_s_2),
	.datab(curr_blk_s_3),
	.datac(curr_blk_s_2),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(cout_1),
	.cout());
defparam \cout[1]~0 .lut_mask = 16'hFFFE;
defparam \cout[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \sum_out[1]~0 (
	.dataa(curr_blk_s_3),
	.datab(addr_s_2),
	.datac(curr_blk_s_2),
	.datad(addr_s_1),
	.cin(gnd),
	.combout(sum_out_1),
	.cout());
defparam \sum_out[1]~0 .lut_mask = 16'h6996;
defparam \sum_out[1]~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_core (
	curr_blk_s_1,
	curr_blk_s_0,
	Add0,
	Add01,
	out_stall_d,
	curr_pwr_2_s,
	out_valid,
	enable,
	out_enable,
	processing,
	processing1,
	out_valid1,
	cnt_1,
	cnt_0,
	cnt_2,
	in_eop,
	out_real_0,
	out_real_1,
	out_real_2,
	out_real_3,
	out_real_4,
	out_real_5,
	out_real_6,
	out_real_7,
	out_imag_0,
	out_imag_1,
	out_imag_2,
	out_imag_3,
	out_imag_4,
	out_imag_5,
	out_imag_6,
	out_imag_7,
	out_data_8,
	out_data_0,
	curr_inverse_s,
	out_data_9,
	out_data_1,
	out_data_10,
	out_data_2,
	out_data_11,
	out_data_3,
	out_data_12,
	out_data_4,
	out_data_13,
	out_data_5,
	out_data_14,
	out_data_6,
	out_data_15,
	out_data_7,
	curr_input_sel_s_0,
	Add02,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_1;
input 	curr_blk_s_0;
input 	Add0;
input 	Add01;
input 	out_stall_d;
input 	curr_pwr_2_s;
output 	out_valid;
input 	enable;
output 	out_enable;
output 	processing;
output 	processing1;
output 	out_valid1;
input 	cnt_1;
input 	cnt_0;
input 	cnt_2;
input 	in_eop;
output 	out_real_0;
output 	out_real_1;
output 	out_real_2;
output 	out_real_3;
output 	out_real_4;
output 	out_real_5;
output 	out_real_6;
output 	out_real_7;
output 	out_imag_0;
output 	out_imag_1;
output 	out_imag_2;
output 	out_imag_3;
output 	out_imag_4;
output 	out_imag_5;
output 	out_imag_6;
output 	out_imag_7;
input 	out_data_8;
input 	out_data_0;
input 	curr_inverse_s;
input 	out_data_9;
input 	out_data_1;
input 	out_data_10;
input 	out_data_2;
input 	out_data_11;
input 	out_data_3;
input 	out_data_12;
input 	out_data_4;
input 	out_data_13;
input 	out_data_5;
input 	out_data_14;
input 	out_data_6;
input 	out_data_15;
input 	out_data_7;
input 	curr_input_sel_s_0;
input 	Add02;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~0_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[2]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~0_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[2]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~1_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[3]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~1_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[3]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~2_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[4]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~2_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[4]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~3_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[5]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~3_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[5]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~4_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[6]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~4_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[6]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~5_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[7]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~5_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[7]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~6_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[8]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~6_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[8]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~7_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[9]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~7_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[9]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[0]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[1]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[2]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[3]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[4]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[5]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[6]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[7]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[2]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ;
wire \ena_ctrl|sop~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_valid~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_inverse_next~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[9]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[9]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_inverse~q ;
wire \stg_in_sop[0]~0_combout ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_eop~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_sop_next~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_eop_next~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_sop~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[0]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[1]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[2]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[3]~q ;
wire \gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[1]~q ;
wire \stg_in_imag[0][2]~0_combout ;
wire \stg_in_imag[0][1]~1_combout ;
wire \stg_in_imag[0][0]~2_combout ;
wire \stg_in_real[0][2]~0_combout ;
wire \stg_in_real[0][1]~1_combout ;
wire \stg_in_real[0][0]~2_combout ;
wire \stg_in_imag[0][3]~3_combout ;
wire \stg_in_real[0][3]~3_combout ;
wire \stg_in_imag[0][4]~4_combout ;
wire \stg_in_real[0][4]~4_combout ;
wire \stg_in_imag[0][5]~5_combout ;
wire \stg_in_real[0][5]~5_combout ;
wire \stg_in_imag[0][6]~6_combout ;
wire \stg_in_real[0][6]~6_combout ;
wire \stg_in_imag[0][7]~7_combout ;
wire \stg_in_real[0][7]~7_combout ;
wire \stg_in_sop[0]~1_combout ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[0]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[1]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[2]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[3]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[4]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[5]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[6]~q ;
wire \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[7]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[1]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[2]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[0]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[1]~q ;
wire \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[2]~q ;
wire \gen_natural_order_core:gen_stages:1:r22_stage|twid_rd_en~0_combout ;
wire \out_imag[0]~0_combout ;
wire \out_imag[0]~1_combout ;
wire \out_inverse~0_combout ;
wire \out_imag[1]~2_combout ;
wire \out_imag[1]~3_combout ;
wire \out_imag[2]~4_combout ;
wire \out_imag[2]~5_combout ;
wire \out_imag[3]~6_combout ;
wire \out_imag[3]~7_combout ;
wire \out_imag[4]~8_combout ;
wire \out_imag[4]~9_combout ;
wire \out_imag[5]~10_combout ;
wire \out_imag[5]~11_combout ;
wire \out_imag[6]~12_combout ;
wire \out_imag[6]~13_combout ;
wire \out_imag[7]~14_combout ;
wire \out_imag[7]~15_combout ;


ifft_8p_auk_dspip_r22sdf_twrom \gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2 (
	.imagtwid_0(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[0]~q ),
	.imagtwid_1(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[1]~q ),
	.imagtwid_2(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[2]~q ),
	.imagtwid_3(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[3]~q ),
	.imagtwid_4(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[4]~q ),
	.imagtwid_5(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[5]~q ),
	.imagtwid_6(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[6]~q ),
	.imagtwid_7(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[7]~q ),
	.curr_blk_s_1(curr_blk_s_1),
	.stg_valid_next(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ),
	.curr_pwr_2_s(curr_pwr_2_s),
	.enable(out_enable),
	.realtwid_0(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[0]~q ),
	.realtwid_1(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[1]~q ),
	.realtwid_2(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[2]~q ),
	.realtwid_3(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[3]~q ),
	.realtwid_4(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[4]~q ),
	.realtwid_5(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[5]~q ),
	.realtwid_6(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[6]~q ),
	.realtwid_7(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[7]~q ),
	.control_s_1(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[1]~q ),
	.control_s_2(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[2]~q ),
	.control_s_0(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[0]~q ),
	.rd_en(\gen_natural_order_core:gen_stages:1:r22_stage|twid_rd_en~0_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset(reset_n));

ifft_8p_auk_dspip_r22sdf_stage_1 \gen_natural_order_core:gen_stages:1:r22_stage (
	.stg_imag_next_0(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~q ),
	.stg_real_next_0(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~q ),
	.stg_imag_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~q ),
	.stg_real_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~q ),
	.stg_imag_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~q ),
	.stg_real_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~q ),
	.stg_imag_next_3(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~q ),
	.stg_real_next_3(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~q ),
	.stg_imag_next_4(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~q ),
	.stg_real_next_4(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~q ),
	.stg_imag_next_5(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~q ),
	.stg_real_next_5(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~q ),
	.stg_imag_next_6(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~q ),
	.stg_real_next_6(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~q ),
	.stg_imag_next_7(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~q ),
	.stg_real_next_7(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~q ),
	.imagtwid_0(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[0]~q ),
	.imagtwid_1(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[1]~q ),
	.imagtwid_2(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[2]~q ),
	.imagtwid_3(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[3]~q ),
	.imagtwid_4(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[4]~q ),
	.imagtwid_5(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[5]~q ),
	.imagtwid_6(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[6]~q ),
	.imagtwid_7(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|imagtwid[7]~q ),
	.curr_blk_s_1(curr_blk_s_1),
	.out_stall_d(out_stall_d),
	.out_valid(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ),
	.stg_valid_next(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(\ena_ctrl|sop~q ),
	.out_valid_s(enable),
	.out_enable(out_enable),
	.processing1(processing1),
	.out_imag_2(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ),
	.out_real_2(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ),
	.out_inverse(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ),
	.stg_inverse_next(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_inverse_next~q ),
	.out_imag_3(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ),
	.out_real_3(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ),
	.out_imag_4(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ),
	.out_real_4(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ),
	.out_imag_5(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ),
	.out_real_5(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ),
	.out_imag_6(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ),
	.out_real_6(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ),
	.out_imag_7(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ),
	.out_real_7(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ),
	.out_imag_8(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ),
	.out_real_8(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ),
	.out_imag_9(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[9]~q ),
	.out_real_9(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[9]~q ),
	.stg_sop_next(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_sop_next~q ),
	.stg_eop_next(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_eop_next~q ),
	.fftpts_less_one_0(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[0]~q ),
	.fftpts_less_one_1(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[1]~q ),
	.fftpts_less_one_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[2]~q ),
	.fftpts_less_one_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[3]~q ),
	.realtwid_0(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[0]~q ),
	.realtwid_1(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[1]~q ),
	.realtwid_2(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[2]~q ),
	.realtwid_3(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[3]~q ),
	.realtwid_4(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[4]~q ),
	.realtwid_5(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[5]~q ),
	.realtwid_6(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[6]~q ),
	.realtwid_7(\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|realtwid[7]~q ),
	.control_s_1(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[1]~q ),
	.control_s_2(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[2]~q ),
	.control_s_0(\gen_natural_order_core:gen_stages:1:r22_stage|gen_cma:cma_inst|bf_counter_inst|control_s[0]~q ),
	.stg_control_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[1]~q ),
	.stg_control_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[2]~q ),
	.twid_rd_en(\gen_natural_order_core:gen_stages:1:r22_stage|twid_rd_en~0_combout ),
	.clk(clk),
	.reset(reset_n));

ifft_8p_auk_dspip_r22sdf_stg_pipe \gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect (
	.stg_imag_next_0(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~q ),
	.stg_real_next_0(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~q ),
	.stg_imag_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~q ),
	.stg_real_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~q ),
	.stg_imag_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~q ),
	.stg_real_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~q ),
	.stg_imag_next_3(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~q ),
	.stg_real_next_3(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~q ),
	.stg_imag_next_4(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~q ),
	.stg_real_next_4(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~q ),
	.stg_imag_next_5(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~q ),
	.stg_real_next_5(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~q ),
	.stg_imag_next_6(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~q ),
	.stg_real_next_6(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~q ),
	.stg_imag_next_7(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~q ),
	.stg_real_next_7(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~q ),
	.stg_imag_next_01(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~0_combout ),
	.out_imag_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[2]~q ),
	.stg_real_next_01(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~0_combout ),
	.out_real_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[2]~q ),
	.stg_imag_next_11(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~1_combout ),
	.out_imag_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[3]~q ),
	.stg_real_next_11(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~1_combout ),
	.out_real_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[3]~q ),
	.stg_imag_next_21(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~2_combout ),
	.out_imag_4(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[4]~q ),
	.stg_real_next_21(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~2_combout ),
	.out_real_4(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[4]~q ),
	.stg_imag_next_31(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~3_combout ),
	.out_imag_5(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[5]~q ),
	.stg_real_next_31(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~3_combout ),
	.out_real_5(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[5]~q ),
	.stg_imag_next_41(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~4_combout ),
	.out_imag_6(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[6]~q ),
	.stg_real_next_41(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~4_combout ),
	.out_real_6(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[6]~q ),
	.stg_imag_next_51(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~5_combout ),
	.out_imag_7(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[7]~q ),
	.stg_real_next_51(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~5_combout ),
	.out_real_7(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[7]~q ),
	.stg_imag_next_61(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~6_combout ),
	.out_imag_8(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[8]~q ),
	.stg_real_next_61(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~6_combout ),
	.out_real_8(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[8]~q ),
	.stg_imag_next_71(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~7_combout ),
	.out_imag_9(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[9]~q ),
	.stg_real_next_71(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~7_combout ),
	.out_real_9(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[9]~q ),
	.out_control_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[2]~q ),
	.curr_blk_s_1(curr_blk_s_1),
	.stg_valid_next1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ),
	.out_valid_s(enable),
	.out_enable(out_enable),
	.out_valid(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_valid~q ),
	.Equal1(in_eop),
	.stg_inverse_next1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_inverse_next~q ),
	.out_data_8(out_data_8),
	.out_data_0(out_data_0),
	.curr_inverse_s(curr_inverse_s),
	.out_inverse(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_inverse~q ),
	.out_data_9(out_data_9),
	.out_data_1(out_data_1),
	.out_data_10(out_data_10),
	.out_data_2(out_data_2),
	.out_data_11(out_data_11),
	.out_data_3(out_data_3),
	.out_data_12(out_data_12),
	.out_data_4(out_data_4),
	.out_data_13(out_data_13),
	.out_data_5(out_data_5),
	.out_data_14(out_data_14),
	.out_data_6(out_data_6),
	.out_data_15(out_data_15),
	.out_data_7(out_data_7),
	.stg_in_sop_0(\stg_in_sop[0]~0_combout ),
	.out_eop(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_eop~q ),
	.stg_sop_next1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_sop_next~q ),
	.stg_eop_next1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_eop_next~q ),
	.out_sop(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_sop~q ),
	.out_control_1(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[1]~q ),
	.stg_control_next_1(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[1]~q ),
	.stg_control_next_2(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_control_next[2]~q ),
	.clk(clk),
	.reset_n(reset_n));

ifft_8p_auk_dspip_r22sdf_stage \gen_natural_order_core:gen_stages:0:r22_stage (
	.out_imag_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[2]~q ),
	.out_real_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[2]~q ),
	.out_imag_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[3]~q ),
	.out_real_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[3]~q ),
	.out_imag_4(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[4]~q ),
	.out_real_4(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[4]~q ),
	.out_imag_5(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[5]~q ),
	.out_real_5(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[5]~q ),
	.out_imag_6(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[6]~q ),
	.out_real_6(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[6]~q ),
	.out_imag_7(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[7]~q ),
	.out_real_7(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[7]~q ),
	.out_imag_8(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[8]~q ),
	.out_real_8(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[8]~q ),
	.out_imag_9(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_imag[9]~q ),
	.out_real_9(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_real[9]~q ),
	.out_control_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[2]~q ),
	.curr_blk_s_0(curr_blk_s_0),
	.Add0(Add0),
	.Add01(Add01),
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(\ena_ctrl|sop~q ),
	.out_valid_s(enable),
	.out_enable(out_enable),
	.processing1(processing),
	.out_valid(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_valid~q ),
	.curr_inverse_s(curr_inverse_s),
	.out_inverse(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_inverse~q ),
	.curr_input_sel_s_0(curr_input_sel_s_0),
	.stg_in_sop_0(\stg_in_sop[0]~0_combout ),
	.out_eop(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_eop~q ),
	.out_sop(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|out_sop~q ),
	.fftpts_less_one_0(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[0]~q ),
	.fftpts_less_one_1(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[1]~q ),
	.fftpts_less_one_2(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[2]~q ),
	.fftpts_less_one_3(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|bf_control_inst|fftpts_less_one[3]~q ),
	.Add02(Add02),
	.out_control_1(\gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|bf_control_inst|out_control[1]~q ),
	.stg_in_imag_2_0(\stg_in_imag[0][2]~0_combout ),
	.stg_in_imag_1_0(\stg_in_imag[0][1]~1_combout ),
	.stg_in_imag_0_0(\stg_in_imag[0][0]~2_combout ),
	.stg_in_real_2_0(\stg_in_real[0][2]~0_combout ),
	.stg_in_real_1_0(\stg_in_real[0][1]~1_combout ),
	.stg_in_real_0_0(\stg_in_real[0][0]~2_combout ),
	.stg_in_imag_3_0(\stg_in_imag[0][3]~3_combout ),
	.stg_in_real_3_0(\stg_in_real[0][3]~3_combout ),
	.stg_in_imag_4_0(\stg_in_imag[0][4]~4_combout ),
	.stg_in_real_4_0(\stg_in_real[0][4]~4_combout ),
	.stg_in_imag_5_0(\stg_in_imag[0][5]~5_combout ),
	.stg_in_real_5_0(\stg_in_real[0][5]~5_combout ),
	.stg_in_imag_6_0(\stg_in_imag[0][6]~6_combout ),
	.stg_in_real_6_0(\stg_in_real[0][6]~6_combout ),
	.stg_in_imag_7_0(\stg_in_imag[0][7]~7_combout ),
	.stg_in_real_7_0(\stg_in_real[0][7]~7_combout ),
	.stg_in_sop_01(\stg_in_sop[0]~1_combout ),
	.clk(clk),
	.reset(reset_n));

ifft_8p_auk_dspip_r22sdf_enable_control ena_ctrl(
	.out_stall_d(out_stall_d),
	.sop1(\ena_ctrl|sop~q ),
	.enable(enable),
	.out_enable(out_enable),
	.in_eop(in_eop),
	.clk(clk),
	.reset_n(reset_n));

cycloneiv_lcell_comb \stg_in_sop[0]~0 (
	.dataa(gnd),
	.datab(cnt_2),
	.datac(cnt_0),
	.datad(cnt_1),
	.cin(gnd),
	.combout(\stg_in_sop[0]~0_combout ),
	.cout());
defparam \stg_in_sop[0]~0 .lut_mask = 16'h3FFF;
defparam \stg_in_sop[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][2]~0 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~2_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][2]~0_combout ),
	.cout());
defparam \stg_in_imag[0][2]~0 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][2]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][1]~1 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~1_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][1]~1_combout ),
	.cout());
defparam \stg_in_imag[0][1]~1 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][0]~2 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~0_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][0]~2_combout ),
	.cout());
defparam \stg_in_imag[0][0]~2 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][0]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][2]~0 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~2_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][2]~0_combout ),
	.cout());
defparam \stg_in_real[0][2]~0 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][2]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][1]~1 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~1_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][1]~1_combout ),
	.cout());
defparam \stg_in_real[0][1]~1 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][0]~2 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~0_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][0]~2_combout ),
	.cout());
defparam \stg_in_real[0][0]~2 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][0]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][3]~3 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~3_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][3]~3_combout ),
	.cout());
defparam \stg_in_imag[0][3]~3 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][3]~3 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~3_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][3]~3_combout ),
	.cout());
defparam \stg_in_real[0][3]~3 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][4]~4 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~4_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][4]~4_combout ),
	.cout());
defparam \stg_in_imag[0][4]~4 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][4]~4 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~4_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][4]~4_combout ),
	.cout());
defparam \stg_in_real[0][4]~4 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][5]~5 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~5_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][5]~5_combout ),
	.cout());
defparam \stg_in_imag[0][5]~5 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][5]~5 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~5_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][5]~5_combout ),
	.cout());
defparam \stg_in_real[0][5]~5 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][6]~6 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~6_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][6]~6_combout ),
	.cout());
defparam \stg_in_imag[0][6]~6 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][6]~6 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~6_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][6]~6_combout ),
	.cout());
defparam \stg_in_real[0][6]~6 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_imag[0][7]~7 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~7_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_imag[0][7]~7_combout ),
	.cout());
defparam \stg_in_imag[0][7]~7 .lut_mask = 16'hEEEE;
defparam \stg_in_imag[0][7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_real[0][7]~7 (
	.dataa(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~7_combout ),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\stg_in_real[0][7]~7_combout ),
	.cout());
defparam \stg_in_real[0][7]~7 .lut_mask = 16'hEEEE;
defparam \stg_in_real[0][7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_in_sop[0]~1 (
	.dataa(curr_input_sel_s_0),
	.datab(cnt_2),
	.datac(cnt_0),
	.datad(cnt_1),
	.cin(gnd),
	.combout(\stg_in_sop[0]~1_combout ),
	.cout());
defparam \stg_in_sop[0]~1 .lut_mask = 16'hBFFF;
defparam \stg_in_sop[0]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_valid~0 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(out_valid),
	.cout());
defparam \out_valid~0 .lut_mask = 16'hAACC;
defparam \out_valid~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_valid~1 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_valid_next~q ),
	.datac(curr_pwr_2_s),
	.datad(out_enable),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam \out_valid~1 .lut_mask = 16'hFFAC;
defparam \out_valid~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[0]~0 (
	.dataa(\out_imag[0]~0_combout ),
	.datab(\out_imag[0]~1_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_0),
	.cout());
defparam \out_real[0]~0 .lut_mask = 16'hAACC;
defparam \out_real[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[1]~1 (
	.dataa(\out_imag[1]~2_combout ),
	.datab(\out_imag[1]~3_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_1),
	.cout());
defparam \out_real[1]~1 .lut_mask = 16'hAACC;
defparam \out_real[1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[2]~2 (
	.dataa(\out_imag[2]~4_combout ),
	.datab(\out_imag[2]~5_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_2),
	.cout());
defparam \out_real[2]~2 .lut_mask = 16'hAACC;
defparam \out_real[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[3]~3 (
	.dataa(\out_imag[3]~6_combout ),
	.datab(\out_imag[3]~7_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_3),
	.cout());
defparam \out_real[3]~3 .lut_mask = 16'hAACC;
defparam \out_real[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[4]~4 (
	.dataa(\out_imag[4]~8_combout ),
	.datab(\out_imag[4]~9_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_4),
	.cout());
defparam \out_real[4]~4 .lut_mask = 16'hAACC;
defparam \out_real[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[5]~5 (
	.dataa(\out_imag[5]~10_combout ),
	.datab(\out_imag[5]~11_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_5),
	.cout());
defparam \out_real[5]~5 .lut_mask = 16'hAACC;
defparam \out_real[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[6]~6 (
	.dataa(\out_imag[6]~12_combout ),
	.datab(\out_imag[6]~13_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_6),
	.cout());
defparam \out_real[6]~6 .lut_mask = 16'hAACC;
defparam \out_real[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_real[7]~7 (
	.dataa(\out_imag[7]~14_combout ),
	.datab(\out_imag[7]~15_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_real_7),
	.cout());
defparam \out_real[7]~7 .lut_mask = 16'hAACC;
defparam \out_real[7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[0]~16 (
	.dataa(\out_imag[0]~1_combout ),
	.datab(\out_imag[0]~0_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_0),
	.cout());
defparam \out_imag[0]~16 .lut_mask = 16'hAACC;
defparam \out_imag[0]~16 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[1]~17 (
	.dataa(\out_imag[1]~3_combout ),
	.datab(\out_imag[1]~2_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_1),
	.cout());
defparam \out_imag[1]~17 .lut_mask = 16'hAACC;
defparam \out_imag[1]~17 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[2]~18 (
	.dataa(\out_imag[2]~5_combout ),
	.datab(\out_imag[2]~4_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_2),
	.cout());
defparam \out_imag[2]~18 .lut_mask = 16'hAACC;
defparam \out_imag[2]~18 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[3]~19 (
	.dataa(\out_imag[3]~7_combout ),
	.datab(\out_imag[3]~6_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_3),
	.cout());
defparam \out_imag[3]~19 .lut_mask = 16'hAACC;
defparam \out_imag[3]~19 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[4]~20 (
	.dataa(\out_imag[4]~9_combout ),
	.datab(\out_imag[4]~8_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_4),
	.cout());
defparam \out_imag[4]~20 .lut_mask = 16'hAACC;
defparam \out_imag[4]~20 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[5]~21 (
	.dataa(\out_imag[5]~11_combout ),
	.datab(\out_imag[5]~10_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_5),
	.cout());
defparam \out_imag[5]~21 .lut_mask = 16'hAACC;
defparam \out_imag[5]~21 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[6]~22 (
	.dataa(\out_imag[6]~13_combout ),
	.datab(\out_imag[6]~12_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_6),
	.cout());
defparam \out_imag[6]~22 .lut_mask = 16'hAACC;
defparam \out_imag[6]~22 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[7]~23 (
	.dataa(\out_imag[7]~15_combout ),
	.datab(\out_imag[7]~14_combout ),
	.datac(gnd),
	.datad(\out_inverse~0_combout ),
	.cin(gnd),
	.combout(out_imag_7),
	.cout());
defparam \out_imag[7]~23 .lut_mask = 16'hAACC;
defparam \out_imag[7]~23 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[0]~0 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[0]~0_combout ),
	.cout());
defparam \out_imag[0]~0 .lut_mask = 16'hAACC;
defparam \out_imag[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[0]~1 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[0]~1_combout ),
	.cout());
defparam \out_imag[0]~1 .lut_mask = 16'hAACC;
defparam \out_imag[0]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_inverse~0 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_inverse_next~q ),
	.datac(curr_pwr_2_s),
	.datad(out_enable),
	.cin(gnd),
	.combout(\out_inverse~0_combout ),
	.cout());
defparam \out_inverse~0 .lut_mask = 16'hFFAC;
defparam \out_inverse~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[1]~2 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[1]~2_combout ),
	.cout());
defparam \out_imag[1]~2 .lut_mask = 16'hAACC;
defparam \out_imag[1]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[1]~3 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[1]~3_combout ),
	.cout());
defparam \out_imag[1]~3 .lut_mask = 16'hAACC;
defparam \out_imag[1]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[2]~4 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[2]~4_combout ),
	.cout());
defparam \out_imag[2]~4 .lut_mask = 16'hAACC;
defparam \out_imag[2]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[2]~5 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[2]~5_combout ),
	.cout());
defparam \out_imag[2]~5 .lut_mask = 16'hAACC;
defparam \out_imag[2]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[3]~6 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[3]~6_combout ),
	.cout());
defparam \out_imag[3]~6 .lut_mask = 16'hAACC;
defparam \out_imag[3]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[3]~7 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[3]~7_combout ),
	.cout());
defparam \out_imag[3]~7 .lut_mask = 16'hAACC;
defparam \out_imag[3]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[4]~8 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[4]~8_combout ),
	.cout());
defparam \out_imag[4]~8 .lut_mask = 16'hAACC;
defparam \out_imag[4]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[4]~9 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[4]~9_combout ),
	.cout());
defparam \out_imag[4]~9 .lut_mask = 16'hAACC;
defparam \out_imag[4]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[5]~10 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[5]~10_combout ),
	.cout());
defparam \out_imag[5]~10 .lut_mask = 16'hAACC;
defparam \out_imag[5]~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[5]~11 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[5]~11_combout ),
	.cout());
defparam \out_imag[5]~11 .lut_mask = 16'hAACC;
defparam \out_imag[5]~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[6]~12 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[6]~12_combout ),
	.cout());
defparam \out_imag[6]~12 .lut_mask = 16'hAACC;
defparam \out_imag[6]~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[6]~13 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[6]~13_combout ),
	.cout());
defparam \out_imag[6]~13 .lut_mask = 16'hAACC;
defparam \out_imag[6]~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[7]~14 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_imag[9]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_imag_next[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[7]~14_combout ),
	.cout());
defparam \out_imag[7]~14 .lut_mask = 16'hAACC;
defparam \out_imag[7]~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_imag[7]~15 (
	.dataa(\gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|out_real[9]~q ),
	.datab(\gen_natural_order_core:gen_stages:0:gen_stg_connect:stg_connect|stg_real_next[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag[7]~15_combout ),
	.cout());
defparam \out_imag[7]~15 .lut_mask = 16'hAACC;
defparam \out_imag[7]~15 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_enable_control (
	out_stall_d,
	sop1,
	enable,
	out_enable,
	in_eop,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
input 	out_stall_d;
output 	sop1;
input 	enable;
output 	out_enable;
input 	in_eop;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



dffeas sop(
	.clk(clk),
	.d(in_eop),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(sop1),
	.prn(vcc));
defparam sop.is_wysiwyg = "true";
defparam sop.power_up = "low";

cycloneiv_lcell_comb \out_enable~0 (
	.dataa(out_stall_d),
	.datab(gnd),
	.datac(sop1),
	.datad(enable),
	.cin(gnd),
	.combout(out_enable),
	.cout());
defparam \out_enable~0 .lut_mask = 16'hF505;
defparam \out_enable~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_stage (
	out_imag_2,
	out_real_2,
	out_imag_3,
	out_real_3,
	out_imag_4,
	out_real_4,
	out_imag_5,
	out_real_5,
	out_imag_6,
	out_real_6,
	out_imag_7,
	out_real_7,
	out_imag_8,
	out_real_8,
	out_imag_9,
	out_real_9,
	out_control_2,
	curr_blk_s_0,
	Add0,
	Add01,
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	out_enable,
	processing1,
	out_valid,
	curr_inverse_s,
	out_inverse,
	curr_input_sel_s_0,
	stg_in_sop_0,
	out_eop,
	out_sop,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	Add02,
	out_control_1,
	stg_in_imag_2_0,
	stg_in_imag_1_0,
	stg_in_imag_0_0,
	stg_in_real_2_0,
	stg_in_real_1_0,
	stg_in_real_0_0,
	stg_in_imag_3_0,
	stg_in_real_3_0,
	stg_in_imag_4_0,
	stg_in_real_4_0,
	stg_in_imag_5_0,
	stg_in_real_5_0,
	stg_in_imag_6_0,
	stg_in_real_6_0,
	stg_in_imag_7_0,
	stg_in_real_7_0,
	stg_in_sop_01,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	out_imag_2;
output 	out_real_2;
output 	out_imag_3;
output 	out_real_3;
output 	out_imag_4;
output 	out_real_4;
output 	out_imag_5;
output 	out_real_5;
output 	out_imag_6;
output 	out_real_6;
output 	out_imag_7;
output 	out_real_7;
output 	out_imag_8;
output 	out_real_8;
output 	out_imag_9;
output 	out_real_9;
output 	out_control_2;
input 	curr_blk_s_0;
input 	Add0;
input 	Add01;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	out_enable;
output 	processing1;
output 	out_valid;
input 	curr_inverse_s;
output 	out_inverse;
input 	curr_input_sel_s_0;
input 	stg_in_sop_0;
output 	out_eop;
output 	out_sop;
output 	fftpts_less_one_0;
output 	fftpts_less_one_1;
output 	fftpts_less_one_2;
output 	fftpts_less_one_3;
input 	Add02;
output 	out_control_1;
input 	stg_in_imag_2_0;
input 	stg_in_imag_1_0;
input 	stg_in_imag_0_0;
input 	stg_in_real_2_0;
input 	stg_in_real_1_0;
input 	stg_in_real_0_0;
input 	stg_in_imag_3_0;
input 	stg_in_real_3_0;
input 	stg_in_imag_4_0;
input 	stg_in_real_4_0;
input 	stg_in_imag_5_0;
input 	stg_in_real_5_0;
input 	stg_in_imag_6_0;
input 	stg_in_real_6_0;
input 	stg_in_imag_7_0;
input 	stg_in_real_7_0;
input 	stg_in_sop_01;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[1]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[1]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[0]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[0]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_sop~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ;
wire \processing_bfi_cnt_p~0_combout ;
wire \processing_cnt[0]~1_combout ;
wire \processing_cnt[2]~0_combout ;
wire \processing_cnt[0]~q ;
wire \Add2~1_combout ;
wire \processing_cnt[1]~q ;
wire \Add2~0_combout ;
wire \processing_cnt[2]~q ;
wire \res~0_combout ;


ifft_8p_auk_dspip_r22sdf_bfii \gen_bfii:bfii_inst (
	.out_imag_2(out_imag_2),
	.out_real_2(out_real_2),
	.out_imag_3(out_imag_3),
	.out_real_3(out_real_3),
	.out_imag_4(out_imag_4),
	.out_real_4(out_real_4),
	.out_imag_5(out_imag_5),
	.out_real_5(out_real_5),
	.out_imag_6(out_imag_6),
	.out_real_6(out_real_6),
	.out_imag_7(out_imag_7),
	.out_real_7(out_real_7),
	.out_imag_8(out_imag_8),
	.out_real_8(out_real_8),
	.out_imag_9(out_imag_9),
	.out_real_9(out_real_9),
	.out_imag_21(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ),
	.out_real_21(\gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ),
	.out_imag_1(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[1]~q ),
	.out_real_1(\gen_bfi:gen_bfi_only:bfi_inst|out_real[1]~q ),
	.out_imag_0(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[0]~q ),
	.out_real_0(\gen_bfi:gen_bfi_only:bfi_inst|out_real[0]~q ),
	.out_imag_31(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ),
	.out_real_31(\gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ),
	.out_imag_41(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ),
	.out_real_41(\gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ),
	.out_imag_51(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ),
	.out_real_51(\gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ),
	.out_imag_61(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ),
	.out_real_61(\gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ),
	.out_imag_71(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ),
	.out_real_71(\gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ),
	.out_imag_81(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ),
	.out_real_81(\gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ),
	.out_control_2(out_control_2),
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(out_enable),
	.out_valid1(out_valid),
	.out_inverse1(out_inverse),
	.out_eop1(out_eop),
	.out_sop1(out_sop),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.out_sop2(\gen_bfi:gen_bfi_only:bfi_inst|out_sop~q ),
	.out_valid2(\gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ),
	.out_inverse2(\gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ),
	.out_control_1(out_control_1),
	.clk(clk),
	.reset(reset));

ifft_8p_auk_dspip_r22sdf_bfi \gen_bfi:gen_bfi_only:bfi_inst (
	.out_imag_2(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[2]~q ),
	.out_real_2(\gen_bfi:gen_bfi_only:bfi_inst|out_real[2]~q ),
	.out_imag_1(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[1]~q ),
	.out_real_1(\gen_bfi:gen_bfi_only:bfi_inst|out_real[1]~q ),
	.out_imag_0(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[0]~q ),
	.out_real_0(\gen_bfi:gen_bfi_only:bfi_inst|out_real[0]~q ),
	.out_imag_3(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[3]~q ),
	.out_real_3(\gen_bfi:gen_bfi_only:bfi_inst|out_real[3]~q ),
	.out_imag_4(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[4]~q ),
	.out_real_4(\gen_bfi:gen_bfi_only:bfi_inst|out_real[4]~q ),
	.out_imag_5(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[5]~q ),
	.out_real_5(\gen_bfi:gen_bfi_only:bfi_inst|out_real[5]~q ),
	.out_imag_6(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[6]~q ),
	.out_real_6(\gen_bfi:gen_bfi_only:bfi_inst|out_real[6]~q ),
	.out_imag_7(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[7]~q ),
	.out_real_7(\gen_bfi:gen_bfi_only:bfi_inst|out_real[7]~q ),
	.out_imag_8(\gen_bfi:gen_bfi_only:bfi_inst|out_imag[8]~q ),
	.out_real_8(\gen_bfi:gen_bfi_only:bfi_inst|out_real[8]~q ),
	.curr_blk_s_0(curr_blk_s_0),
	.Add0(Add0),
	.Add01(Add01),
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(out_enable),
	.curr_inverse_s(curr_inverse_s),
	.curr_input_sel_s_0(curr_input_sel_s_0),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.Add02(Add02),
	.out_sop1(\gen_bfi:gen_bfi_only:bfi_inst|out_sop~q ),
	.out_valid1(\gen_bfi:gen_bfi_only:bfi_inst|out_valid~q ),
	.out_inverse1(\gen_bfi:gen_bfi_only:bfi_inst|out_inverse~q ),
	.in_imag({gnd,stg_in_imag_7_0,stg_in_imag_6_0,stg_in_imag_5_0,stg_in_imag_4_0,stg_in_imag_3_0,stg_in_imag_2_0,stg_in_imag_1_0,stg_in_imag_0_0}),
	.in_real({gnd,stg_in_real_7_0,stg_in_real_6_0,stg_in_real_5_0,stg_in_real_4_0,stg_in_real_3_0,stg_in_real_2_0,stg_in_real_1_0,stg_in_real_0_0}),
	.stg_in_sop_0(stg_in_sop_01),
	.clk(clk),
	.reset(reset));

dffeas processing(
	.clk(clk),
	.d(\res~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(processing1),
	.prn(vcc));
defparam processing.is_wysiwyg = "true";
defparam processing.power_up = "low";

cycloneiv_lcell_comb \processing_bfi_cnt_p~0 (
	.dataa(gnd),
	.datab(out_valid_s),
	.datac(curr_input_sel_s_0),
	.datad(stg_in_sop_0),
	.cin(gnd),
	.combout(\processing_bfi_cnt_p~0_combout ),
	.cout());
defparam \processing_bfi_cnt_p~0 .lut_mask = 16'h3FFF;
defparam \processing_bfi_cnt_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[0]~1 (
	.dataa(\processing_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\processing_cnt[0]~1_combout ),
	.cout());
defparam \processing_cnt[0]~1 .lut_mask = 16'h5555;
defparam \processing_cnt[0]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[2]~0 (
	.dataa(out_enable),
	.datab(\processing_bfi_cnt_p~0_combout ),
	.datac(out_valid),
	.datad(out_eop),
	.cin(gnd),
	.combout(\processing_cnt[2]~0_combout ),
	.cout());
defparam \processing_cnt[2]~0 .lut_mask = 16'hEBBE;
defparam \processing_cnt[2]~0 .sum_lutc_input = "datac";

dffeas \processing_cnt[0] (
	.clk(clk),
	.d(\processing_cnt[0]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~0_combout ),
	.q(\processing_cnt[0]~q ),
	.prn(vcc));
defparam \processing_cnt[0] .is_wysiwyg = "true";
defparam \processing_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \Add2~1 (
	.dataa(\processing_cnt[1]~q ),
	.datab(\processing_cnt[0]~q ),
	.datac(\processing_bfi_cnt_p~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h9696;
defparam \Add2~1 .sum_lutc_input = "datac";

dffeas \processing_cnt[1] (
	.clk(clk),
	.d(\Add2~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~0_combout ),
	.q(\processing_cnt[1]~q ),
	.prn(vcc));
defparam \processing_cnt[1] .is_wysiwyg = "true";
defparam \processing_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Add2~0 (
	.dataa(\processing_cnt[2]~q ),
	.datab(\processing_bfi_cnt_p~0_combout ),
	.datac(\processing_cnt[1]~q ),
	.datad(\processing_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h6996;
defparam \Add2~0 .sum_lutc_input = "datac";

dffeas \processing_cnt[2] (
	.clk(clk),
	.d(\Add2~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~0_combout ),
	.q(\processing_cnt[2]~q ),
	.prn(vcc));
defparam \processing_cnt[2] .is_wysiwyg = "true";
defparam \processing_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \res~0 (
	.dataa(\processing_cnt[2]~q ),
	.datab(\processing_cnt[1]~q ),
	.datac(\processing_cnt[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\res~0_combout ),
	.cout());
defparam \res~0 .lut_mask = 16'hFEFE;
defparam \res~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_bfi (
	out_imag_2,
	out_real_2,
	out_imag_1,
	out_real_1,
	out_imag_0,
	out_real_0,
	out_imag_3,
	out_real_3,
	out_imag_4,
	out_real_4,
	out_imag_5,
	out_real_5,
	out_imag_6,
	out_real_6,
	out_imag_7,
	out_real_7,
	out_imag_8,
	out_real_8,
	curr_blk_s_0,
	Add0,
	Add01,
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	curr_inverse_s,
	curr_input_sel_s_0,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	Add02,
	out_sop1,
	out_valid1,
	out_inverse1,
	in_imag,
	in_real,
	stg_in_sop_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	out_imag_2;
output 	out_real_2;
output 	out_imag_1;
output 	out_real_1;
output 	out_imag_0;
output 	out_real_0;
output 	out_imag_3;
output 	out_real_3;
output 	out_imag_4;
output 	out_real_4;
output 	out_imag_5;
output 	out_real_5;
output 	out_imag_6;
output 	out_real_6;
output 	out_imag_7;
output 	out_real_7;
output 	out_imag_8;
output 	out_real_8;
input 	curr_blk_s_0;
input 	Add0;
input 	Add01;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
input 	curr_inverse_s;
input 	curr_input_sel_s_0;
output 	fftpts_less_one_0;
output 	fftpts_less_one_1;
output 	fftpts_less_one_2;
output 	fftpts_less_one_3;
input 	Add02;
output 	out_sop1;
output 	out_valid1;
output 	out_inverse1;
input 	[8:0] in_imag;
input 	[8:0] in_real;
input 	stg_in_sop_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \bf_control_inst|out_sop~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][2]~q ;
wire \generate_delay_less_pipeline:in_imag_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][1]~q ;
wire \generate_delay_less_pipeline:in_imag_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][0]~q ;
wire \generate_delay_less_pipeline:in_imag_d[0]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][2]~q ;
wire \generate_delay_less_pipeline:in_real_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][1]~q ;
wire \generate_delay_less_pipeline:in_real_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][0]~q ;
wire \generate_delay_less_pipeline:in_real_d[0]~q ;
wire \bf_control_inst|out_inverse~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][3]~q ;
wire \generate_delay_less_pipeline:in_imag_d[3]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][3]~q ;
wire \generate_delay_less_pipeline:in_real_d[3]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][4]~q ;
wire \generate_delay_less_pipeline:in_imag_d[4]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][4]~q ;
wire \generate_delay_less_pipeline:in_real_d[4]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][5]~q ;
wire \generate_delay_less_pipeline:in_imag_d[5]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][5]~q ;
wire \generate_delay_less_pipeline:in_real_d[5]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][6]~q ;
wire \generate_delay_less_pipeline:in_imag_d[6]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][6]~q ;
wire \generate_delay_less_pipeline:in_real_d[6]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[3][7]~q ;
wire \generate_delay_less_pipeline:in_imag_d[7]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[3][7]~q ;
wire \generate_delay_less_pipeline:in_real_d[7]~q ;
wire \bf_control_inst|bf_counter_inst|control_s[2]~q ;
wire \bf_control_inst|out_valid~combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][2]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ;
wire \del_in_imag_pl_d~0_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][1]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ;
wire \del_in_imag_pl_d~1_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][0]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ;
wire \del_in_imag_pl_d~2_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][2]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ;
wire \del_in_real_pl_d~0_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][1]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ;
wire \del_in_real_pl_d~1_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][0]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ;
wire \del_in_real_pl_d~2_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][3]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ;
wire \del_in_imag_pl_d~3_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][3]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ;
wire \del_in_real_pl_d~3_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][4]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ;
wire \del_in_imag_pl_d~4_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][4]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ;
wire \del_in_real_pl_d~4_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][5]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ;
wire \del_in_imag_pl_d~5_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][5]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ;
wire \del_in_real_pl_d~5_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][6]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ;
wire \del_in_imag_pl_d~6_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][6]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ;
wire \del_in_real_pl_d~6_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[2][7]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ;
wire \del_in_imag_pl_d~7_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][7]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ;
wire \del_in_real_pl_d~7_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ;
wire \del_in_imag_pl_d~8_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ;
wire \del_in_imag_pl_d~9_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ;
wire \del_in_imag_pl_d~10_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ;
wire \del_in_real_pl_d~8_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ;
wire \del_in_real_pl_d~9_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ;
wire \del_in_real_pl_d~10_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ;
wire \del_in_imag_pl_d~11_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ;
wire \del_in_real_pl_d~11_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ;
wire \del_in_imag_pl_d~12_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ;
wire \del_in_real_pl_d~12_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ;
wire \del_in_imag_pl_d~13_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ;
wire \del_in_real_pl_d~13_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ;
wire \del_in_imag_pl_d~14_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ;
wire \del_in_real_pl_d~14_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][8]~q ;
wire \del_in_imag_pl_d~15_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][8]~q ;
wire \del_in_real_pl_d~15_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][2]~q ;
wire \out_imag~0_combout ;
wire \s_sel_d[0]~q ;
wire \s_sel_d[1]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][2]~q ;
wire \out_real~0_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][1]~q ;
wire \out_imag~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][1]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][1]~q ;
wire \out_real~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][0]~q ;
wire \out_imag~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][0]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][0]~q ;
wire \out_real~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][3]~q ;
wire \out_imag~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][3]~q ;
wire \out_real~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][4]~q ;
wire \out_imag~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][4]~q ;
wire \out_real~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][5]~q ;
wire \out_imag~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][5]~q ;
wire \out_real~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][6]~q ;
wire \out_imag~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][6]~q ;
wire \out_real~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][7]~q ;
wire \out_imag~7_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][7]~q ;
wire \out_real~7_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[2][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[3][8]~q ;
wire \out_imag~8_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[2][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[3][8]~q ;
wire \out_real~8_combout ;
wire \out_sop_d[0]~q ;
wire \out_valid_d[0]~q ;
wire \out_valid_d[1]~q ;
wire \out_inverse_d[0]~q ;


ifft_8p_auk_dspip_r22sdf_bf_control bf_control_inst(
	.curr_blk_s_0(curr_blk_s_0),
	.Add0(Add0),
	.Add01(Add01),
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(enable),
	.curr_inverse_s(curr_inverse_s),
	.curr_input_sel_s_0(curr_input_sel_s_0),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.Add02(Add02),
	.out_sop1(\bf_control_inst|out_sop~q ),
	.out_inverse1(\bf_control_inst|out_inverse~q ),
	.control_s_2(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.out_valid1(\bf_control_inst|out_valid~combout ),
	.stg_in_sop_0(stg_in_sop_0),
	.clk(clk),
	.reset(reset));

ifft_8p_auk_dspip_r22sdf_addsub_2 \gen_fixedpt_adders:in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(\generate_delay_less_pipeline:del_in_imag_pl_d[3][2]~q ),
	.generate_delay_less_pipelinein_imag_d2(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(\generate_delay_less_pipeline:del_in_imag_pl_d[3][1]~q ),
	.generate_delay_less_pipelinein_imag_d1(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(\generate_delay_less_pipeline:del_in_imag_pl_d[3][0]~q ),
	.generate_delay_less_pipelinein_imag_d0(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(\generate_delay_less_pipeline:del_in_imag_pl_d[3][3]~q ),
	.generate_delay_less_pipelinein_imag_d3(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(\generate_delay_less_pipeline:del_in_imag_pl_d[3][4]~q ),
	.generate_delay_less_pipelinein_imag_d4(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(\generate_delay_less_pipeline:del_in_imag_pl_d[3][5]~q ),
	.generate_delay_less_pipelinein_imag_d5(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(\generate_delay_less_pipeline:del_in_imag_pl_d[3][6]~q ),
	.generate_delay_less_pipelinein_imag_d6(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(\generate_delay_less_pipeline:del_in_imag_pl_d[3][7]~q ),
	.generate_delay_less_pipelinein_imag_d7(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_3 \gen_fixedpt_adders:in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d32(\generate_delay_less_pipeline:del_in_real_pl_d[3][2]~q ),
	.generate_delay_less_pipelinein_real_d2(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d31(\generate_delay_less_pipeline:del_in_real_pl_d[3][1]~q ),
	.generate_delay_less_pipelinein_real_d1(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d30(\generate_delay_less_pipeline:del_in_real_pl_d[3][0]~q ),
	.generate_delay_less_pipelinein_real_d0(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d33(\generate_delay_less_pipeline:del_in_real_pl_d[3][3]~q ),
	.generate_delay_less_pipelinein_real_d3(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d34(\generate_delay_less_pipeline:del_in_real_pl_d[3][4]~q ),
	.generate_delay_less_pipelinein_real_d4(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d35(\generate_delay_less_pipeline:del_in_real_pl_d[3][5]~q ),
	.generate_delay_less_pipelinein_real_d5(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d36(\generate_delay_less_pipeline:del_in_real_pl_d[3][6]~q ),
	.generate_delay_less_pipelinein_real_d6(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d37(\generate_delay_less_pipeline:del_in_real_pl_d[3][7]~q ),
	.generate_delay_less_pipelinein_real_d7(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub \gen_fixedpt_adders:del_in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(\generate_delay_less_pipeline:del_in_imag_pl_d[3][2]~q ),
	.generate_delay_less_pipelinein_imag_d2(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(\generate_delay_less_pipeline:del_in_imag_pl_d[3][1]~q ),
	.generate_delay_less_pipelinein_imag_d1(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(\generate_delay_less_pipeline:del_in_imag_pl_d[3][0]~q ),
	.generate_delay_less_pipelinein_imag_d0(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(\generate_delay_less_pipeline:del_in_imag_pl_d[3][3]~q ),
	.generate_delay_less_pipelinein_imag_d3(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(\generate_delay_less_pipeline:del_in_imag_pl_d[3][4]~q ),
	.generate_delay_less_pipelinein_imag_d4(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(\generate_delay_less_pipeline:del_in_imag_pl_d[3][5]~q ),
	.generate_delay_less_pipelinein_imag_d5(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(\generate_delay_less_pipeline:del_in_imag_pl_d[3][6]~q ),
	.generate_delay_less_pipelinein_imag_d6(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(\generate_delay_less_pipeline:del_in_imag_pl_d[3][7]~q ),
	.generate_delay_less_pipelinein_imag_d7(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_1 \gen_fixedpt_adders:del_in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_1(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.pipeline_dffe_0(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d32(\generate_delay_less_pipeline:del_in_real_pl_d[3][2]~q ),
	.generate_delay_less_pipelinein_real_d2(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d31(\generate_delay_less_pipeline:del_in_real_pl_d[3][1]~q ),
	.generate_delay_less_pipelinein_real_d1(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d30(\generate_delay_less_pipeline:del_in_real_pl_d[3][0]~q ),
	.generate_delay_less_pipelinein_real_d0(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d33(\generate_delay_less_pipeline:del_in_real_pl_d[3][3]~q ),
	.generate_delay_less_pipelinein_real_d3(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d34(\generate_delay_less_pipeline:del_in_real_pl_d[3][4]~q ),
	.generate_delay_less_pipelinein_real_d4(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d35(\generate_delay_less_pipeline:del_in_real_pl_d[3][5]~q ),
	.generate_delay_less_pipelinein_real_d5(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d36(\generate_delay_less_pipeline:del_in_real_pl_d[3][6]~q ),
	.generate_delay_less_pipelinein_real_d6(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d37(\generate_delay_less_pipeline:del_in_real_pl_d[3][7]~q ),
	.generate_delay_less_pipelinein_real_d7(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][2] (
	.clk(clk),
	.d(\del_in_imag_pl_d~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[2] (
	.clk(clk),
	.d(in_imag[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][1] (
	.clk(clk),
	.d(\del_in_imag_pl_d~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[1] (
	.clk(clk),
	.d(in_imag[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][0] (
	.clk(clk),
	.d(\del_in_imag_pl_d~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[0] (
	.clk(clk),
	.d(in_imag[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][2] (
	.clk(clk),
	.d(\del_in_real_pl_d~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[2] (
	.clk(clk),
	.d(in_real[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][1] (
	.clk(clk),
	.d(\del_in_real_pl_d~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[1] (
	.clk(clk),
	.d(in_real[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][0] (
	.clk(clk),
	.d(\del_in_real_pl_d~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[0] (
	.clk(clk),
	.d(in_real[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][3] (
	.clk(clk),
	.d(\del_in_imag_pl_d~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[3] (
	.clk(clk),
	.d(in_imag[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][3] (
	.clk(clk),
	.d(\del_in_real_pl_d~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[3] (
	.clk(clk),
	.d(in_real[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][4] (
	.clk(clk),
	.d(\del_in_imag_pl_d~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[4] (
	.clk(clk),
	.d(in_imag[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][4] (
	.clk(clk),
	.d(\del_in_real_pl_d~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[4] (
	.clk(clk),
	.d(in_real[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][5] (
	.clk(clk),
	.d(\del_in_imag_pl_d~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[5] (
	.clk(clk),
	.d(in_imag[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][5] (
	.clk(clk),
	.d(\del_in_real_pl_d~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[5] (
	.clk(clk),
	.d(in_real[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][6] (
	.clk(clk),
	.d(\del_in_imag_pl_d~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[6] (
	.clk(clk),
	.d(in_imag[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][6] (
	.clk(clk),
	.d(\del_in_real_pl_d~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[6] (
	.clk(clk),
	.d(in_real[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[3][7] (
	.clk(clk),
	.d(\del_in_imag_pl_d~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[3][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[3][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[7] (
	.clk(clk),
	.d(in_imag[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[3][7] (
	.clk(clk),
	.d(\del_in_real_pl_d~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[3][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[3][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[7] (
	.clk(clk),
	.d(in_real[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] (
	.clk(clk),
	.d(\del_in_imag_pl_d~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~0 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][2]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~0_combout ),
	.cout());
defparam \del_in_imag_pl_d~0 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] (
	.clk(clk),
	.d(\del_in_imag_pl_d~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~1 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][1]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~1_combout ),
	.cout());
defparam \del_in_imag_pl_d~1 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] (
	.clk(clk),
	.d(\del_in_imag_pl_d~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~2 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][0]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~2_combout ),
	.cout());
defparam \del_in_imag_pl_d~2 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][2] (
	.clk(clk),
	.d(\del_in_real_pl_d~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~0 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][2]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~0_combout ),
	.cout());
defparam \del_in_real_pl_d~0 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][1] (
	.clk(clk),
	.d(\del_in_real_pl_d~9_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~1 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][1]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~1_combout ),
	.cout());
defparam \del_in_real_pl_d~1 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][0] (
	.clk(clk),
	.d(\del_in_real_pl_d~10_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~2 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][0]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~2_combout ),
	.cout());
defparam \del_in_real_pl_d~2 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] (
	.clk(clk),
	.d(\del_in_imag_pl_d~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~3 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][3]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~3_combout ),
	.cout());
defparam \del_in_imag_pl_d~3 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][3] (
	.clk(clk),
	.d(\del_in_real_pl_d~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~3 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][3]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~3_combout ),
	.cout());
defparam \del_in_real_pl_d~3 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] (
	.clk(clk),
	.d(\del_in_imag_pl_d~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~4 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][4]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~4_combout ),
	.cout());
defparam \del_in_imag_pl_d~4 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][4] (
	.clk(clk),
	.d(\del_in_real_pl_d~12_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~4 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][4]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~4_combout ),
	.cout());
defparam \del_in_real_pl_d~4 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] (
	.clk(clk),
	.d(\del_in_imag_pl_d~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~5 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][5]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~5_combout ),
	.cout());
defparam \del_in_imag_pl_d~5 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][5] (
	.clk(clk),
	.d(\del_in_real_pl_d~13_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~5 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][5]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~5_combout ),
	.cout());
defparam \del_in_real_pl_d~5 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] (
	.clk(clk),
	.d(\del_in_imag_pl_d~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~6 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][6]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~6_combout ),
	.cout());
defparam \del_in_imag_pl_d~6 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][6] (
	.clk(clk),
	.d(\del_in_real_pl_d~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~6 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][6]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~6_combout ),
	.cout());
defparam \del_in_real_pl_d~6 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[2][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[2][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[2][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] (
	.clk(clk),
	.d(\del_in_imag_pl_d~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~7 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[2][7]~q ),
	.datab(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~7_combout ),
	.cout());
defparam \del_in_imag_pl_d~7 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[2][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][7] (
	.clk(clk),
	.d(\del_in_real_pl_d~15_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][7] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~7 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~q ),
	.datab(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~7_combout ),
	.cout());
defparam \del_in_real_pl_d~7 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0 (
	.dataa(curr_pwr_2_s),
	.datab(out_valid_s),
	.datac(sop),
	.datad(out_stall_d),
	.cin(gnd),
	.combout(\generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0_combout ),
	.cout());
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0 .lut_mask = 16'hACFF;
defparam \generate_delay_less_pipeline:del_in_real_pl_d[2][7]~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~8 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~8_combout ),
	.cout());
defparam \del_in_imag_pl_d~8 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~8 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~9 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~9_combout ),
	.cout());
defparam \del_in_imag_pl_d~9 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~9 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~10 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~10_combout ),
	.cout());
defparam \del_in_imag_pl_d~10 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~10 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~8 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~8_combout ),
	.cout());
defparam \del_in_real_pl_d~8 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~8 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~9 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~9_combout ),
	.cout());
defparam \del_in_real_pl_d~9 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~9 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~10 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~10_combout ),
	.cout());
defparam \del_in_real_pl_d~10 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~10 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~11 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~11_combout ),
	.cout());
defparam \del_in_imag_pl_d~11 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~11 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~11 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~11_combout ),
	.cout());
defparam \del_in_real_pl_d~11 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~11 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~12 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~12_combout ),
	.cout());
defparam \del_in_imag_pl_d~12 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~12 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~12 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~12_combout ),
	.cout());
defparam \del_in_real_pl_d~12 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~12 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~13 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~13_combout ),
	.cout());
defparam \del_in_imag_pl_d~13 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~13 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~13 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~13_combout ),
	.cout());
defparam \del_in_real_pl_d~13 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~13 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~14 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~14_combout ),
	.cout());
defparam \del_in_imag_pl_d~14 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~14 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~14 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~14_combout ),
	.cout());
defparam \del_in_real_pl_d~14 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~14 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][8] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~15 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][8]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~15_combout ),
	.cout());
defparam \del_in_imag_pl_d~15 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~15 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][8] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~15 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][8]~q ),
	.datab(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~15_combout ),
	.cout());
defparam \del_in_real_pl_d~15 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~15 .sum_lutc_input = "datac";

dffeas \out_imag[2] (
	.clk(clk),
	.d(\out_imag~0_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_2),
	.prn(vcc));
defparam \out_imag[2] .is_wysiwyg = "true";
defparam \out_imag[2] .power_up = "low";

dffeas \out_real[2] (
	.clk(clk),
	.d(\out_real~0_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_2),
	.prn(vcc));
defparam \out_real[2] .is_wysiwyg = "true";
defparam \out_real[2] .power_up = "low";

dffeas \out_imag[1] (
	.clk(clk),
	.d(\out_imag~1_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_1),
	.prn(vcc));
defparam \out_imag[1] .is_wysiwyg = "true";
defparam \out_imag[1] .power_up = "low";

dffeas \out_real[1] (
	.clk(clk),
	.d(\out_real~1_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_1),
	.prn(vcc));
defparam \out_real[1] .is_wysiwyg = "true";
defparam \out_real[1] .power_up = "low";

dffeas \out_imag[0] (
	.clk(clk),
	.d(\out_imag~2_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_0),
	.prn(vcc));
defparam \out_imag[0] .is_wysiwyg = "true";
defparam \out_imag[0] .power_up = "low";

dffeas \out_real[0] (
	.clk(clk),
	.d(\out_real~2_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_0),
	.prn(vcc));
defparam \out_real[0] .is_wysiwyg = "true";
defparam \out_real[0] .power_up = "low";

dffeas \out_imag[3] (
	.clk(clk),
	.d(\out_imag~3_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_3),
	.prn(vcc));
defparam \out_imag[3] .is_wysiwyg = "true";
defparam \out_imag[3] .power_up = "low";

dffeas \out_real[3] (
	.clk(clk),
	.d(\out_real~3_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_3),
	.prn(vcc));
defparam \out_real[3] .is_wysiwyg = "true";
defparam \out_real[3] .power_up = "low";

dffeas \out_imag[4] (
	.clk(clk),
	.d(\out_imag~4_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_4),
	.prn(vcc));
defparam \out_imag[4] .is_wysiwyg = "true";
defparam \out_imag[4] .power_up = "low";

dffeas \out_real[4] (
	.clk(clk),
	.d(\out_real~4_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_4),
	.prn(vcc));
defparam \out_real[4] .is_wysiwyg = "true";
defparam \out_real[4] .power_up = "low";

dffeas \out_imag[5] (
	.clk(clk),
	.d(\out_imag~5_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_5),
	.prn(vcc));
defparam \out_imag[5] .is_wysiwyg = "true";
defparam \out_imag[5] .power_up = "low";

dffeas \out_real[5] (
	.clk(clk),
	.d(\out_real~5_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_5),
	.prn(vcc));
defparam \out_real[5] .is_wysiwyg = "true";
defparam \out_real[5] .power_up = "low";

dffeas \out_imag[6] (
	.clk(clk),
	.d(\out_imag~6_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_6),
	.prn(vcc));
defparam \out_imag[6] .is_wysiwyg = "true";
defparam \out_imag[6] .power_up = "low";

dffeas \out_real[6] (
	.clk(clk),
	.d(\out_real~6_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_6),
	.prn(vcc));
defparam \out_real[6] .is_wysiwyg = "true";
defparam \out_real[6] .power_up = "low";

dffeas \out_imag[7] (
	.clk(clk),
	.d(\out_imag~7_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_7),
	.prn(vcc));
defparam \out_imag[7] .is_wysiwyg = "true";
defparam \out_imag[7] .power_up = "low";

dffeas \out_real[7] (
	.clk(clk),
	.d(\out_real~7_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_7),
	.prn(vcc));
defparam \out_real[7] .is_wysiwyg = "true";
defparam \out_real[7] .power_up = "low";

dffeas \out_imag[8] (
	.clk(clk),
	.d(\out_imag~8_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_8),
	.prn(vcc));
defparam \out_imag[8] .is_wysiwyg = "true";
defparam \out_imag[8] .power_up = "low";

dffeas \out_real[8] (
	.clk(clk),
	.d(\out_real~8_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_8),
	.prn(vcc));
defparam \out_real[8] .is_wysiwyg = "true";
defparam \out_real[8] .power_up = "low";

dffeas out_sop(
	.clk(clk),
	.d(\out_sop_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_sop1),
	.prn(vcc));
defparam out_sop.is_wysiwyg = "true";
defparam out_sop.power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\out_valid_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][2] .power_up = "low";

cycloneiv_lcell_comb \out_imag~0 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~0_combout ),
	.cout());
defparam \out_imag~0 .lut_mask = 16'hAACC;
defparam \out_imag~0 .sum_lutc_input = "datac";

dffeas \s_sel_d[0] (
	.clk(clk),
	.d(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[0]~q ),
	.prn(vcc));
defparam \s_sel_d[0] .is_wysiwyg = "true";
defparam \s_sel_d[0] .power_up = "low";

dffeas \s_sel_d[1] (
	.clk(clk),
	.d(\s_sel_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[1]~q ),
	.prn(vcc));
defparam \s_sel_d[1] .is_wysiwyg = "true";
defparam \s_sel_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][2] .power_up = "low";

cycloneiv_lcell_comb \out_real~0 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~0_combout ),
	.cout());
defparam \out_real~0 .lut_mask = 16'hAACC;
defparam \out_real~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][1] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][1] .power_up = "low";

cycloneiv_lcell_comb \out_imag~1 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][1]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~1_combout ),
	.cout());
defparam \out_imag~1 .lut_mask = 16'hAACC;
defparam \out_imag~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][1] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][1] .power_up = "low";

cycloneiv_lcell_comb \out_real~1 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][1]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~1_combout ),
	.cout());
defparam \out_real~1 .lut_mask = 16'hAACC;
defparam \out_real~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][0] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][0] .power_up = "low";

cycloneiv_lcell_comb \out_imag~2 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][0]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~2_combout ),
	.cout());
defparam \out_imag~2 .lut_mask = 16'hAACC;
defparam \out_imag~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][0] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][0] .power_up = "low";

cycloneiv_lcell_comb \out_real~2 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][0]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~2_combout ),
	.cout());
defparam \out_real~2 .lut_mask = 16'hAACC;
defparam \out_real~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][3] .power_up = "low";

cycloneiv_lcell_comb \out_imag~3 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~3_combout ),
	.cout());
defparam \out_imag~3 .lut_mask = 16'hAACC;
defparam \out_imag~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][3] .power_up = "low";

cycloneiv_lcell_comb \out_real~3 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~3_combout ),
	.cout());
defparam \out_real~3 .lut_mask = 16'hAACC;
defparam \out_real~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][4] .power_up = "low";

cycloneiv_lcell_comb \out_imag~4 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~4_combout ),
	.cout());
defparam \out_imag~4 .lut_mask = 16'hAACC;
defparam \out_imag~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][4] .power_up = "low";

cycloneiv_lcell_comb \out_real~4 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~4_combout ),
	.cout());
defparam \out_real~4 .lut_mask = 16'hAACC;
defparam \out_real~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][5] .power_up = "low";

cycloneiv_lcell_comb \out_imag~5 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~5_combout ),
	.cout());
defparam \out_imag~5 .lut_mask = 16'hAACC;
defparam \out_imag~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][5] .power_up = "low";

cycloneiv_lcell_comb \out_real~5 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~5_combout ),
	.cout());
defparam \out_real~5 .lut_mask = 16'hAACC;
defparam \out_real~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][6] .power_up = "low";

cycloneiv_lcell_comb \out_imag~6 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~6_combout ),
	.cout());
defparam \out_imag~6 .lut_mask = 16'hAACC;
defparam \out_imag~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][6] .power_up = "low";

cycloneiv_lcell_comb \out_real~6 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~6_combout ),
	.cout());
defparam \out_real~6 .lut_mask = 16'hAACC;
defparam \out_real~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][7] .power_up = "low";

cycloneiv_lcell_comb \out_imag~7 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~7_combout ),
	.cout());
defparam \out_imag~7 .lut_mask = 16'hAACC;
defparam \out_imag~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][7] .power_up = "low";

cycloneiv_lcell_comb \out_real~7 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~7_combout ),
	.cout());
defparam \out_real~7 .lut_mask = 16'hAACC;
defparam \out_real~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[2][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[2][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[2][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[3][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[2][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[3][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[3][8] .power_up = "low";

cycloneiv_lcell_comb \out_imag~8 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[3][8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~8_combout ),
	.cout());
defparam \out_imag~8 .lut_mask = 16'hAACC;
defparam \out_imag~8 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[2][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[2][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[2][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[3][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[2][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[3][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[3][8] .power_up = "low";

cycloneiv_lcell_comb \out_real~8 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[3][8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~8_combout ),
	.cout());
defparam \out_real~8 .lut_mask = 16'hAACC;
defparam \out_real~8 .sum_lutc_input = "datac";

dffeas \out_sop_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_sop~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_sop_d[0]~q ),
	.prn(vcc));
defparam \out_sop_d[0] .is_wysiwyg = "true";
defparam \out_sop_d[0] .power_up = "low";

dffeas \out_valid_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_valid~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[0]~q ),
	.prn(vcc));
defparam \out_valid_d[0] .is_wysiwyg = "true";
defparam \out_valid_d[0] .power_up = "low";

dffeas \out_valid_d[1] (
	.clk(clk),
	.d(\out_valid_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[1]~q ),
	.prn(vcc));
defparam \out_valid_d[1] .is_wysiwyg = "true";
defparam \out_valid_d[1] .power_up = "low";

dffeas \out_inverse_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_inverse~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_inverse_d[0]~q ),
	.prn(vcc));
defparam \out_inverse_d[0] .is_wysiwyg = "true";
defparam \out_inverse_d[0] .power_up = "low";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	out_enable,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_1 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_1 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_sgj auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_sgj (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.datab(generate_delay_less_pipelinein_imag_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .lut_mask = 16'h66EE;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.datab(generate_delay_less_pipelinein_imag_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.datab(generate_delay_less_pipelinein_imag_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.datab(generate_delay_less_pipelinein_imag_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.datab(generate_delay_less_pipelinein_imag_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.datab(generate_delay_less_pipelinein_imag_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.datab(generate_delay_less_pipelinein_imag_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_1 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_2 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d32(generate_delay_less_pipelinedel_in_real_pl_d32),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d31(generate_delay_less_pipelinedel_in_real_pl_d31),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d30(generate_delay_less_pipelinedel_in_real_pl_d30),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d33(generate_delay_less_pipelinedel_in_real_pl_d33),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d34(generate_delay_less_pipelinedel_in_real_pl_d34),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d35(generate_delay_less_pipelinedel_in_real_pl_d35),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d36(generate_delay_less_pipelinedel_in_real_pl_d36),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d37(generate_delay_less_pipelinedel_in_real_pl_d37),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_2 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_sgj_1 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d32(generate_delay_less_pipelinedel_in_real_pl_d32),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d31(generate_delay_less_pipelinedel_in_real_pl_d31),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d30(generate_delay_less_pipelinedel_in_real_pl_d30),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d33(generate_delay_less_pipelinedel_in_real_pl_d33),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d34(generate_delay_less_pipelinedel_in_real_pl_d34),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d35(generate_delay_less_pipelinedel_in_real_pl_d35),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d36(generate_delay_less_pipelinedel_in_real_pl_d36),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d37(generate_delay_less_pipelinedel_in_real_pl_d37),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_sgj_1 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d30),
	.datab(generate_delay_less_pipelinein_real_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .lut_mask = 16'h66EE;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d31),
	.datab(generate_delay_less_pipelinein_real_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d32),
	.datab(generate_delay_less_pipelinein_real_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d33),
	.datab(generate_delay_less_pipelinein_real_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d34),
	.datab(generate_delay_less_pipelinein_real_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d35),
	.datab(generate_delay_less_pipelinein_real_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d36),
	.datab(generate_delay_less_pipelinein_real_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d37),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d37),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_2 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	out_enable,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_3 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_3 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_sgj_2 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_imag_pl_d32(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d31(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d30(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d33(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d34(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d35(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d36(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d37(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_sgj_2 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d32,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d31,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d30,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d33,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d34,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d35,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d36,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d37,
	generate_delay_less_pipelinein_imag_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d32;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d31;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d30;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d33;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d34;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d35;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d36;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d37;
input 	generate_delay_less_pipelinein_imag_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d30),
	.datab(generate_delay_less_pipelinein_imag_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .lut_mask = 16'h66BB;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d31),
	.datab(generate_delay_less_pipelinein_imag_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d32),
	.datab(generate_delay_less_pipelinein_imag_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d33),
	.datab(generate_delay_less_pipelinein_imag_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d34),
	.datab(generate_delay_less_pipelinein_imag_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d35),
	.datab(generate_delay_less_pipelinein_imag_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d36),
	.datab(generate_delay_less_pipelinein_imag_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d37),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_3 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_4 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d32(generate_delay_less_pipelinedel_in_real_pl_d32),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d31(generate_delay_less_pipelinedel_in_real_pl_d31),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d30(generate_delay_less_pipelinedel_in_real_pl_d30),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d33(generate_delay_less_pipelinedel_in_real_pl_d33),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d34(generate_delay_less_pipelinedel_in_real_pl_d34),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d35(generate_delay_less_pipelinedel_in_real_pl_d35),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d36(generate_delay_less_pipelinedel_in_real_pl_d36),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d37(generate_delay_less_pipelinedel_in_real_pl_d37),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_4 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_sgj_3 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_1(pipeline_dffe_1),
	.pipeline_dffe_0(pipeline_dffe_0),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d32(generate_delay_less_pipelinedel_in_real_pl_d32),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d31(generate_delay_less_pipelinedel_in_real_pl_d31),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d30(generate_delay_less_pipelinedel_in_real_pl_d30),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d33(generate_delay_less_pipelinedel_in_real_pl_d33),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d34(generate_delay_less_pipelinedel_in_real_pl_d34),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d35(generate_delay_less_pipelinedel_in_real_pl_d35),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d36(generate_delay_less_pipelinedel_in_real_pl_d36),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d37(generate_delay_less_pipelinedel_in_real_pl_d37),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_sgj_3 (
	pipeline_dffe_2,
	pipeline_dffe_1,
	pipeline_dffe_0,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d32,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d31,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d30,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d33,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d34,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d35,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d36,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d37,
	generate_delay_less_pipelinein_real_d7,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_1;
output 	pipeline_dffe_0;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d32;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d31;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d30;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d33;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d34;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d35;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d36;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d37;
input 	generate_delay_less_pipelinein_real_d7;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_1),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_0),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d30),
	.datab(generate_delay_less_pipelinein_real_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .lut_mask = 16'h66BB;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d31),
	.datab(generate_delay_less_pipelinein_real_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[0]~10 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d32),
	.datab(generate_delay_less_pipelinein_real_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[1]~12 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d33),
	.datab(generate_delay_less_pipelinein_real_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d34),
	.datab(generate_delay_less_pipelinein_real_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d35),
	.datab(generate_delay_less_pipelinein_real_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d36),
	.datab(generate_delay_less_pipelinein_real_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d37),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d37),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_bf_control (
	curr_blk_s_0,
	Add0,
	Add01,
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	curr_inverse_s,
	curr_input_sel_s_0,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	Add02,
	out_sop1,
	out_inverse1,
	control_s_2,
	out_valid1,
	stg_in_sop_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	curr_blk_s_0;
input 	Add0;
input 	Add01;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
input 	curr_inverse_s;
input 	curr_input_sel_s_0;
output 	fftpts_less_one_0;
output 	fftpts_less_one_1;
output 	fftpts_less_one_2;
output 	fftpts_less_one_3;
input 	Add02;
output 	out_sop1;
output 	out_inverse1;
output 	control_s_2;
output 	out_valid1;
input 	stg_in_sop_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fftpts_less_one[0]~0_combout ;
wire \Add3~1_combout ;
wire \in_cnt~3_combout ;
wire \in_cnt[3]~1_combout ;
wire \in_cnt[3]~q ;
wire \Equal0~1_combout ;
wire \in_cnt~2_combout ;
wire \in_cnt[1]~q ;
wire \Equal0~0_combout ;
wire \in_cnt~4_combout ;
wire \in_cnt[0]~q ;
wire \Add3~0_combout ;
wire \in_cnt~0_combout ;
wire \in_cnt[2]~q ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \out_inverse~0_combout ;
wire \out_inverse~1_combout ;
wire \out_cnt[3]~2_combout ;
wire \out_cnt[0]~4_combout ;
wire \out_cnt[0]~q ;
wire \Add4~1_combout ;
wire \out_cnt[2]~6_combout ;
wire \out_cnt[2]~q ;
wire \Add4~0_combout ;
wire \out_cnt[3]~5_combout ;
wire \out_cnt[3]~q ;
wire \out_cnt[0]~0_combout ;
wire \out_cnt[3]~1_combout ;
wire \out_cnt[1]~3_combout ;
wire \out_cnt[1]~q ;
wire \Equal2~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~2_combout ;
wire \shift~4_combout ;
wire \shift~q ;


ifft_8p_auk_dspip_r22sdf_counter bf_counter_inst(
	.curr_pwr_2_s(curr_pwr_2_s),
	.control_s_2(control_s_2),
	.in_cnt_3(\in_cnt[3]~1_combout ),
	.stg_in_sop_0(stg_in_sop_0),
	.clk(clk),
	.reset(reset));

dffeas \fftpts_less_one[0] (
	.clk(clk),
	.d(\fftpts_less_one[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(fftpts_less_one_0),
	.prn(vcc));
defparam \fftpts_less_one[0] .is_wysiwyg = "true";
defparam \fftpts_less_one[0] .power_up = "low";

dffeas \fftpts_less_one[1] (
	.clk(clk),
	.d(Add02),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(fftpts_less_one_1),
	.prn(vcc));
defparam \fftpts_less_one[1] .is_wysiwyg = "true";
defparam \fftpts_less_one[1] .power_up = "low";

dffeas \fftpts_less_one[2] (
	.clk(clk),
	.d(Add01),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(fftpts_less_one_2),
	.prn(vcc));
defparam \fftpts_less_one[2] .is_wysiwyg = "true";
defparam \fftpts_less_one[2] .power_up = "low";

dffeas \fftpts_less_one[3] (
	.clk(clk),
	.d(Add0),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(fftpts_less_one_3),
	.prn(vcc));
defparam \fftpts_less_one[3] .is_wysiwyg = "true";
defparam \fftpts_less_one[3] .power_up = "low";

dffeas out_sop(
	.clk(clk),
	.d(\Equal1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_sop1),
	.prn(vcc));
defparam out_sop.is_wysiwyg = "true";
defparam out_sop.power_up = "low";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

cycloneiv_lcell_comb out_valid(
	.dataa(\shift~q ),
	.datab(control_s_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'hEEEE;
defparam out_valid.sum_lutc_input = "datac";

cycloneiv_lcell_comb \fftpts_less_one[0]~0 (
	.dataa(curr_blk_s_0),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\fftpts_less_one[0]~0_combout ),
	.cout());
defparam \fftpts_less_one[0]~0 .lut_mask = 16'h5555;
defparam \fftpts_less_one[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add3~1 (
	.dataa(\in_cnt[3]~q ),
	.datab(\in_cnt[0]~q ),
	.datac(\in_cnt[1]~q ),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'h6996;
defparam \Add3~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~3 (
	.dataa(\Add3~1_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~3_combout ),
	.cout());
defparam \in_cnt~3 .lut_mask = 16'hAFFF;
defparam \in_cnt~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt[3]~1 (
	.dataa(out_valid_s),
	.datab(curr_input_sel_s_0),
	.datac(sop),
	.datad(out_stall_d),
	.cin(gnd),
	.combout(\in_cnt[3]~1_combout ),
	.cout());
defparam \in_cnt[3]~1 .lut_mask = 16'hFEFF;
defparam \in_cnt[3]~1 .sum_lutc_input = "datac";

dffeas \in_cnt[3] (
	.clk(clk),
	.d(\in_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_cnt[3]~1_combout ),
	.q(\in_cnt[3]~q ),
	.prn(vcc));
defparam \in_cnt[3] .is_wysiwyg = "true";
defparam \in_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \Equal0~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\in_cnt[3]~q ),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~2 (
	.dataa(\in_cnt[0]~q ),
	.datab(\in_cnt[1]~q ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~2_combout ),
	.cout());
defparam \in_cnt~2 .lut_mask = 16'h6FFF;
defparam \in_cnt~2 .sum_lutc_input = "datac";

dffeas \in_cnt[1] (
	.clk(clk),
	.d(\in_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_cnt[3]~1_combout ),
	.q(\in_cnt[1]~q ),
	.prn(vcc));
defparam \in_cnt[1] .is_wysiwyg = "true";
defparam \in_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\in_cnt[1]~q ),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~4 (
	.dataa(\in_cnt[0]~q ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_cnt~4_combout ),
	.cout());
defparam \in_cnt~4 .lut_mask = 16'h7F7F;
defparam \in_cnt~4 .sum_lutc_input = "datac";

dffeas \in_cnt[0] (
	.clk(clk),
	.d(\in_cnt~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_cnt[3]~1_combout ),
	.q(\in_cnt[0]~q ),
	.prn(vcc));
defparam \in_cnt[0] .is_wysiwyg = "true";
defparam \in_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \Add3~0 (
	.dataa(gnd),
	.datab(\in_cnt[2]~q ),
	.datac(\in_cnt[0]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'hC33C;
defparam \Add3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~0 (
	.dataa(\Add3~0_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~0_combout ),
	.cout());
defparam \in_cnt~0 .lut_mask = 16'hAFFF;
defparam \in_cnt~0 .sum_lutc_input = "datac";

dffeas \in_cnt[2] (
	.clk(clk),
	.d(\in_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\in_cnt[3]~1_combout ),
	.q(\in_cnt[2]~q ),
	.prn(vcc));
defparam \in_cnt[2] .is_wysiwyg = "true";
defparam \in_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Equal1~0 (
	.dataa(curr_pwr_2_s),
	.datab(\in_cnt[2]~q ),
	.datac(\in_cnt[1]~q ),
	.datad(\in_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h96FF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal1~1 (
	.dataa(\Equal1~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hAAFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_inverse~0 (
	.dataa(curr_inverse_s),
	.datab(curr_input_sel_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse~0_combout ),
	.cout());
defparam \out_inverse~0 .lut_mask = 16'hEEEE;
defparam \out_inverse~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_inverse~1 (
	.dataa(out_inverse1),
	.datab(\out_inverse~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(enable),
	.cin(gnd),
	.combout(\out_inverse~1_combout ),
	.cout());
defparam \out_inverse~1 .lut_mask = 16'hEFFE;
defparam \out_inverse~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~2 (
	.dataa(\Equal1~1_combout ),
	.datab(\Equal2~2_combout ),
	.datac(\out_cnt[0]~0_combout ),
	.datad(enable),
	.cin(gnd),
	.combout(\out_cnt[3]~2_combout ),
	.cout());
defparam \out_cnt[3]~2 .lut_mask = 16'hFFBF;
defparam \out_cnt[3]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[0]~4 (
	.dataa(\out_cnt[3]~1_combout ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(gnd),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\out_cnt[0]~4_combout ),
	.cout());
defparam \out_cnt[0]~4 .lut_mask = 16'hAACC;
defparam \out_cnt[0]~4 .sum_lutc_input = "datac";

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(\out_cnt[2]~q ),
	.datac(\out_cnt[0]~q ),
	.datad(\out_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add4~1_combout ),
	.cout());
defparam \Add4~1 .lut_mask = 16'hC33C;
defparam \Add4~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[2]~6 (
	.dataa(\out_cnt[2]~q ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(\Add4~1_combout ),
	.datad(\out_cnt[3]~1_combout ),
	.cin(gnd),
	.combout(\out_cnt[2]~6_combout ),
	.cout());
defparam \out_cnt[2]~6 .lut_mask = 16'hFFFE;
defparam \out_cnt[2]~6 .sum_lutc_input = "datac";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Add4~0 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[0]~q ),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout());
defparam \Add4~0 .lut_mask = 16'h6996;
defparam \Add4~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~5 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(\Add4~0_combout ),
	.datad(\out_cnt[3]~1_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~5_combout ),
	.cout());
defparam \out_cnt[3]~5 .lut_mask = 16'hFFFE;
defparam \out_cnt[3]~5 .sum_lutc_input = "datac";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \out_cnt[0]~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\out_cnt[0]~0_combout ),
	.cout());
defparam \out_cnt[0]~0 .lut_mask = 16'h7FFF;
defparam \out_cnt[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~1 (
	.dataa(enable),
	.datab(\out_cnt[0]~0_combout ),
	.datac(\Equal1~1_combout ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~1_combout ),
	.cout());
defparam \out_cnt[3]~1 .lut_mask = 16'hDFFF;
defparam \out_cnt[3]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[1]~3 (
	.dataa(\out_cnt[3]~1_combout ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\out_cnt[1]~3_combout ),
	.cout());
defparam \out_cnt[1]~3 .lut_mask = 16'hEFFE;
defparam \out_cnt[1]~3 .sum_lutc_input = "datac";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal2~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h6996;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal2~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\out_cnt[3]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'h6996;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal2~2 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hEEEE;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shift~4 (
	.dataa(\Equal1~0_combout ),
	.datab(\in_cnt[0]~q ),
	.datac(\shift~q ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(\shift~4_combout ),
	.cout());
defparam \shift~4 .lut_mask = 16'hFBFF;
defparam \shift~4 .sum_lutc_input = "datac";

dffeas shift(
	.clk(clk),
	.d(\shift~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\shift~q ),
	.prn(vcc));
defparam shift.is_wysiwyg = "true";
defparam shift.power_up = "low";

endmodule

module ifft_8p_auk_dspip_r22sdf_counter (
	curr_pwr_2_s,
	control_s_2,
	in_cnt_3,
	stg_in_sop_0,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	curr_pwr_2_s;
output 	control_s_2;
input 	in_cnt_3;
input 	stg_in_sop_0;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_s~2_combout ;
wire \control_s[0]~q ;
wire \control_s~3_combout ;
wire \control_s[1]~q ;
wire \control_s~0_combout ;
wire \control_s~1_combout ;


dffeas \control_s[2] (
	.clk(clk),
	.d(\control_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_cnt_3),
	.q(control_s_2),
	.prn(vcc));
defparam \control_s[2] .is_wysiwyg = "true";
defparam \control_s[2] .power_up = "low";

cycloneiv_lcell_comb \control_s~2 (
	.dataa(curr_pwr_2_s),
	.datab(stg_in_sop_0),
	.datac(gnd),
	.datad(\control_s[0]~q ),
	.cin(gnd),
	.combout(\control_s~2_combout ),
	.cout());
defparam \control_s~2 .lut_mask = 16'h9966;
defparam \control_s~2 .sum_lutc_input = "datac";

dffeas \control_s[0] (
	.clk(clk),
	.d(\control_s~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_cnt_3),
	.q(\control_s[0]~q ),
	.prn(vcc));
defparam \control_s[0] .is_wysiwyg = "true";
defparam \control_s[0] .power_up = "low";

cycloneiv_lcell_comb \control_s~3 (
	.dataa(\control_s[0]~q ),
	.datab(\control_s[1]~q ),
	.datac(stg_in_sop_0),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\control_s~3_combout ),
	.cout());
defparam \control_s~3 .lut_mask = 16'h6996;
defparam \control_s~3 .sum_lutc_input = "datac";

dffeas \control_s[1] (
	.clk(clk),
	.d(\control_s~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(in_cnt_3),
	.q(\control_s[1]~q ),
	.prn(vcc));
defparam \control_s[1] .is_wysiwyg = "true";
defparam \control_s[1] .power_up = "low";

cycloneiv_lcell_comb \control_s~0 (
	.dataa(curr_pwr_2_s),
	.datab(\control_s[0]~q ),
	.datac(control_s_2),
	.datad(\control_s[1]~q ),
	.cin(gnd),
	.combout(\control_s~0_combout ),
	.cout());
defparam \control_s~0 .lut_mask = 16'h6996;
defparam \control_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~1 (
	.dataa(\control_s~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(stg_in_sop_0),
	.cin(gnd),
	.combout(\control_s~1_combout ),
	.cout());
defparam \control_s~1 .lut_mask = 16'hAAFF;
defparam \control_s~1 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_bfii (
	out_imag_2,
	out_real_2,
	out_imag_3,
	out_real_3,
	out_imag_4,
	out_real_4,
	out_imag_5,
	out_real_5,
	out_imag_6,
	out_real_6,
	out_imag_7,
	out_real_7,
	out_imag_8,
	out_real_8,
	out_imag_9,
	out_real_9,
	out_imag_21,
	out_real_21,
	out_imag_1,
	out_real_1,
	out_imag_0,
	out_real_0,
	out_imag_31,
	out_real_31,
	out_imag_41,
	out_real_41,
	out_imag_51,
	out_real_51,
	out_imag_61,
	out_real_61,
	out_imag_71,
	out_real_71,
	out_imag_81,
	out_real_81,
	out_control_2,
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	out_valid1,
	out_inverse1,
	out_eop1,
	out_sop1,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	out_sop2,
	out_valid2,
	out_inverse2,
	out_control_1,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	out_imag_2;
output 	out_real_2;
output 	out_imag_3;
output 	out_real_3;
output 	out_imag_4;
output 	out_real_4;
output 	out_imag_5;
output 	out_real_5;
output 	out_imag_6;
output 	out_real_6;
output 	out_imag_7;
output 	out_real_7;
output 	out_imag_8;
output 	out_real_8;
output 	out_imag_9;
output 	out_real_9;
input 	out_imag_21;
input 	out_real_21;
input 	out_imag_1;
input 	out_real_1;
input 	out_imag_0;
input 	out_real_0;
input 	out_imag_31;
input 	out_real_31;
input 	out_imag_41;
input 	out_real_41;
input 	out_imag_51;
input 	out_real_51;
input 	out_imag_61;
input 	out_real_61;
input 	out_imag_71;
input 	out_real_71;
input 	out_imag_81;
input 	out_real_81;
output 	out_control_2;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
output 	out_valid1;
output 	out_inverse1;
output 	out_eop1;
output 	out_sop1;
input 	fftpts_less_one_0;
input 	fftpts_less_one_1;
input 	fftpts_less_one_2;
input 	fftpts_less_one_3;
input 	out_sop2;
input 	out_valid2;
input 	out_inverse2;
output 	out_control_1;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \bf_control_inst|bf_counter_inst|control_s[1]~q ;
wire \bf_control_inst|out_valid~combout ;
wire \t_sel_d~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[0]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[0]~q ;
wire \bf_control_inst|out_inverse~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[3]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[3]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[4]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[4]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[5]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[5]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[6]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[6]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[7]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[7]~q ;
wire \generate_delay_less_pipeline:in_imag_cmm_d[8]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[1][8]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[1][8]~q ;
wire \generate_delay_less_pipeline:in_real_cmm_d[8]~q ;
wire \bf_control_inst|out_eop~q ;
wire \cmm_control_d~q ;
wire \bf_control_inst|bf_counter_inst|control_s[2]~q ;
wire \in_imag_cmm[2]~0_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ;
wire \del_in_imag_pl_d~0_combout ;
wire \in_imag_cmm[1]~1_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ;
wire \del_in_imag_pl_d~1_combout ;
wire \in_imag_cmm[0]~2_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ;
wire \del_in_imag_pl_d~2_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ;
wire \del_in_real_pl_d~0_combout ;
wire \in_real_cmm[2]~0_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ;
wire \del_in_real_pl_d~1_combout ;
wire \in_real_cmm[1]~1_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ;
wire \del_in_real_pl_d~2_combout ;
wire \in_real_cmm[0]~2_combout ;
wire \in_imag_cmm[3]~3_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ;
wire \del_in_imag_pl_d~3_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ;
wire \del_in_real_pl_d~3_combout ;
wire \in_real_cmm[3]~3_combout ;
wire \in_imag_cmm[4]~4_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ;
wire \del_in_imag_pl_d~4_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ;
wire \del_in_real_pl_d~4_combout ;
wire \in_real_cmm[4]~4_combout ;
wire \in_imag_cmm[5]~5_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ;
wire \del_in_imag_pl_d~5_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ;
wire \del_in_real_pl_d~5_combout ;
wire \in_real_cmm[5]~5_combout ;
wire \in_imag_cmm[6]~6_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ;
wire \del_in_imag_pl_d~6_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ;
wire \del_in_real_pl_d~6_combout ;
wire \in_real_cmm[6]~6_combout ;
wire \in_imag_cmm[7]~7_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ;
wire \del_in_imag_pl_d~7_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ;
wire \del_in_real_pl_d~7_combout ;
wire \in_real_cmm[7]~7_combout ;
wire \in_imag_cmm[8]~8_combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ;
wire \del_in_imag_pl_d~8_combout ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ;
wire \del_in_real_pl_d~8_combout ;
wire \in_real_cmm[8]~8_combout ;
wire \bf_control_inst|out_sop~q ;
wire \cmm_control~combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ;
wire \out_imag~0_combout ;
wire \s_sel_d[0]~q ;
wire \s_sel_d[1]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ;
wire \out_real~0_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ;
wire \out_imag~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ;
wire \out_real~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ;
wire \out_imag~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ;
wire \out_real~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ;
wire \out_imag~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ;
wire \out_real~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ;
wire \out_imag~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ;
wire \out_real~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ;
wire \out_imag~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ;
wire \out_real~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ;
wire \out_imag~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ;
wire \out_real~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[1][9]~q ;
wire \out_imag~7_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ;
wire \generate_delay_less_pipeline:adder2_out_real_d[1][9]~q ;
wire \out_real~7_combout ;
wire \out_valid_d[0]~q ;
wire \out_valid_d[1]~q ;
wire \out_inverse_d[0]~q ;
wire \out_eop_d[0]~q ;
wire \out_sop_d[0]~q ;


ifft_8p_auk_dspip_r22sdf_bf_control_1 bf_control_inst(
	.out_control_2(out_control_2),
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(enable),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.control_s_1(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.out_valid1(\bf_control_inst|out_valid~combout ),
	.out_inverse1(\bf_control_inst|out_inverse~q ),
	.out_eop1(\bf_control_inst|out_eop~q ),
	.out_sop1(out_sop2),
	.out_valid2(out_valid2),
	.control_s_2(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.out_inverse2(out_inverse2),
	.out_sop2(\bf_control_inst|out_sop~q ),
	.out_control_1(out_control_1),
	.clk(clk),
	.reset(reset));

ifft_8p_auk_dspip_r22sdf_addsub_6 \gen_fixedpt_adders:in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinein_imag_cmm_d2(\generate_delay_less_pipeline:in_imag_cmm_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d1(\generate_delay_less_pipeline:in_imag_cmm_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d0(\generate_delay_less_pipeline:in_imag_cmm_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d3(\generate_delay_less_pipeline:in_imag_cmm_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d4(\generate_delay_less_pipeline:in_imag_cmm_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d5(\generate_delay_less_pipeline:in_imag_cmm_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d6(\generate_delay_less_pipeline:in_imag_cmm_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d7(\generate_delay_less_pipeline:in_imag_cmm_d[7]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d8(\generate_delay_less_pipeline:in_imag_cmm_d[8]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(\generate_delay_less_pipeline:del_in_imag_pl_d[1][8]~q ),
	.cmm_control_d(\cmm_control_d~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_7 \gen_fixedpt_adders:in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d12(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.generate_delay_less_pipelinein_real_cmm_d2(\generate_delay_less_pipeline:in_real_cmm_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d11(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.generate_delay_less_pipelinein_real_cmm_d1(\generate_delay_less_pipeline:in_real_cmm_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d10(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.generate_delay_less_pipelinein_real_cmm_d0(\generate_delay_less_pipeline:in_real_cmm_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d13(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.generate_delay_less_pipelinein_real_cmm_d3(\generate_delay_less_pipeline:in_real_cmm_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d14(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.generate_delay_less_pipelinein_real_cmm_d4(\generate_delay_less_pipeline:in_real_cmm_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d15(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.generate_delay_less_pipelinein_real_cmm_d5(\generate_delay_less_pipeline:in_real_cmm_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d16(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.generate_delay_less_pipelinein_real_cmm_d6(\generate_delay_less_pipeline:in_real_cmm_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d17(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.generate_delay_less_pipelinein_real_cmm_d7(\generate_delay_less_pipeline:in_real_cmm_d[7]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d18(\generate_delay_less_pipeline:del_in_real_pl_d[1][8]~q ),
	.generate_delay_less_pipelinein_real_cmm_d8(\generate_delay_less_pipeline:in_real_cmm_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_4 \gen_fixedpt_adders:del_in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.t_sel_d(\t_sel_d~q ),
	.generate_delay_less_pipelinein_imag_cmm_d2(\generate_delay_less_pipeline:in_imag_cmm_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d1(\generate_delay_less_pipeline:in_imag_cmm_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d0(\generate_delay_less_pipeline:in_imag_cmm_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d3(\generate_delay_less_pipeline:in_imag_cmm_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d4(\generate_delay_less_pipeline:in_imag_cmm_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d5(\generate_delay_less_pipeline:in_imag_cmm_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d6(\generate_delay_less_pipeline:in_imag_cmm_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d7(\generate_delay_less_pipeline:in_imag_cmm_d[7]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.generate_delay_less_pipelinein_imag_cmm_d8(\generate_delay_less_pipeline:in_imag_cmm_d[8]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(\generate_delay_less_pipeline:del_in_imag_pl_d[1][8]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_5 \gen_fixedpt_adders:del_in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d12(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.generate_delay_less_pipelinein_real_cmm_d2(\generate_delay_less_pipeline:in_real_cmm_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d11(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.generate_delay_less_pipelinein_real_cmm_d1(\generate_delay_less_pipeline:in_real_cmm_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d10(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.generate_delay_less_pipelinein_real_cmm_d0(\generate_delay_less_pipeline:in_real_cmm_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d13(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.generate_delay_less_pipelinein_real_cmm_d3(\generate_delay_less_pipeline:in_real_cmm_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d14(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.generate_delay_less_pipelinein_real_cmm_d4(\generate_delay_less_pipeline:in_real_cmm_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d15(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.generate_delay_less_pipelinein_real_cmm_d5(\generate_delay_less_pipeline:in_real_cmm_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d16(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.generate_delay_less_pipelinein_real_cmm_d6(\generate_delay_less_pipeline:in_real_cmm_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d17(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.generate_delay_less_pipelinein_real_cmm_d7(\generate_delay_less_pipeline:in_real_cmm_d[7]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d18(\generate_delay_less_pipeline:del_in_real_pl_d[1][8]~q ),
	.generate_delay_less_pipelinein_real_cmm_d8(\generate_delay_less_pipeline:in_real_cmm_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

dffeas t_sel_d(
	.clk(clk),
	.d(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\t_sel_d~q ),
	.prn(vcc));
defparam t_sel_d.is_wysiwyg = "true";
defparam t_sel_d.power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[2] (
	.clk(clk),
	.d(\in_imag_cmm[2]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] (
	.clk(clk),
	.d(\del_in_imag_pl_d~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[1] (
	.clk(clk),
	.d(\in_imag_cmm[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] (
	.clk(clk),
	.d(\del_in_imag_pl_d~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[0] (
	.clk(clk),
	.d(\in_imag_cmm[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] (
	.clk(clk),
	.d(\del_in_imag_pl_d~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][2] (
	.clk(clk),
	.d(\del_in_real_pl_d~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[2] (
	.clk(clk),
	.d(\in_real_cmm[2]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][1] (
	.clk(clk),
	.d(\del_in_real_pl_d~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[1] (
	.clk(clk),
	.d(\in_real_cmm[1]~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][0] (
	.clk(clk),
	.d(\del_in_real_pl_d~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[0] (
	.clk(clk),
	.d(\in_real_cmm[0]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[3] (
	.clk(clk),
	.d(\in_imag_cmm[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] (
	.clk(clk),
	.d(\del_in_imag_pl_d~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][3] (
	.clk(clk),
	.d(\del_in_real_pl_d~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[3] (
	.clk(clk),
	.d(\in_real_cmm[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[4] (
	.clk(clk),
	.d(\in_imag_cmm[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] (
	.clk(clk),
	.d(\del_in_imag_pl_d~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][4] (
	.clk(clk),
	.d(\del_in_real_pl_d~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[4] (
	.clk(clk),
	.d(\in_real_cmm[4]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[5] (
	.clk(clk),
	.d(\in_imag_cmm[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] (
	.clk(clk),
	.d(\del_in_imag_pl_d~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][5] (
	.clk(clk),
	.d(\del_in_real_pl_d~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[5] (
	.clk(clk),
	.d(\in_real_cmm[5]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[6] (
	.clk(clk),
	.d(\in_imag_cmm[6]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] (
	.clk(clk),
	.d(\del_in_imag_pl_d~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][6] (
	.clk(clk),
	.d(\del_in_real_pl_d~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[6] (
	.clk(clk),
	.d(\in_real_cmm[6]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[7] (
	.clk(clk),
	.d(\in_imag_cmm[7]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] (
	.clk(clk),
	.d(\del_in_imag_pl_d~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][7] (
	.clk(clk),
	.d(\del_in_real_pl_d~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[7] (
	.clk(clk),
	.d(\in_real_cmm[7]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_cmm_d[8] (
	.clk(clk),
	.d(\in_imag_cmm[8]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_cmm_d[8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_cmm_d[8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_cmm_d[8] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[1][8] (
	.clk(clk),
	.d(\del_in_imag_pl_d~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[1][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[1][8] (
	.clk(clk),
	.d(\del_in_real_pl_d~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[1][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_cmm_d[8] (
	.clk(clk),
	.d(\in_real_cmm[8]~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_cmm_d[8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_cmm_d[8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_cmm_d[8] .power_up = "low";

dffeas cmm_control_d(
	.clk(clk),
	.d(\cmm_control~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\cmm_control_d~q ),
	.prn(vcc));
defparam cmm_control_d.is_wysiwyg = "true";
defparam cmm_control_d.power_up = "low";

cycloneiv_lcell_comb \in_imag_cmm[2]~0 (
	.dataa(out_imag_21),
	.datab(out_real_21),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[2]~0_combout ),
	.cout());
defparam \in_imag_cmm[2]~0 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[2]~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~0 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~0_combout ),
	.cout());
defparam \del_in_imag_pl_d~0 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[1]~1 (
	.dataa(out_imag_1),
	.datab(out_real_1),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[1]~1_combout ),
	.cout());
defparam \in_imag_cmm[1]~1 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[1]~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~1 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~1_combout ),
	.cout());
defparam \del_in_imag_pl_d~1 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[0]~2 (
	.dataa(out_imag_0),
	.datab(out_real_0),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[0]~2_combout ),
	.cout());
defparam \in_imag_cmm[0]~2 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[0]~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~2 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~2_combout ),
	.cout());
defparam \del_in_imag_pl_d~2 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~0 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~0_combout ),
	.cout());
defparam \del_in_real_pl_d~0 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[2]~0 (
	.dataa(out_real_21),
	.datab(out_imag_21),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[2]~0_combout ),
	.cout());
defparam \in_real_cmm[2]~0 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[2]~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~1 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[1]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~1_combout ),
	.cout());
defparam \del_in_real_pl_d~1 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[1]~1 (
	.dataa(out_real_1),
	.datab(out_imag_1),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[1]~1_combout ),
	.cout());
defparam \in_real_cmm[1]~1 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[1]~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~2 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[0]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~2_combout ),
	.cout());
defparam \del_in_real_pl_d~2 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[0]~2 (
	.dataa(out_real_0),
	.datab(out_imag_0),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[0]~2_combout ),
	.cout());
defparam \in_real_cmm[0]~2 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[0]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[3]~3 (
	.dataa(out_imag_31),
	.datab(out_real_31),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[3]~3_combout ),
	.cout());
defparam \in_imag_cmm[3]~3 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[3]~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~3 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~3_combout ),
	.cout());
defparam \del_in_imag_pl_d~3 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~3 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~3_combout ),
	.cout());
defparam \del_in_real_pl_d~3 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[3]~3 (
	.dataa(out_real_31),
	.datab(out_imag_31),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[3]~3_combout ),
	.cout());
defparam \in_real_cmm[3]~3 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[4]~4 (
	.dataa(out_imag_41),
	.datab(out_real_41),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[4]~4_combout ),
	.cout());
defparam \in_imag_cmm[4]~4 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[4]~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~4 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~4_combout ),
	.cout());
defparam \del_in_imag_pl_d~4 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~4 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~4_combout ),
	.cout());
defparam \del_in_real_pl_d~4 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[4]~4 (
	.dataa(out_real_41),
	.datab(out_imag_41),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[4]~4_combout ),
	.cout());
defparam \in_real_cmm[4]~4 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[5]~5 (
	.dataa(out_imag_51),
	.datab(out_real_51),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[5]~5_combout ),
	.cout());
defparam \in_imag_cmm[5]~5 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[5]~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~5 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~5_combout ),
	.cout());
defparam \del_in_imag_pl_d~5 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~5 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~5_combout ),
	.cout());
defparam \del_in_real_pl_d~5 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[5]~5 (
	.dataa(out_real_51),
	.datab(out_imag_51),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[5]~5_combout ),
	.cout());
defparam \in_real_cmm[5]~5 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[6]~6 (
	.dataa(out_imag_61),
	.datab(out_real_61),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[6]~6_combout ),
	.cout());
defparam \in_imag_cmm[6]~6 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[6]~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~6 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~6_combout ),
	.cout());
defparam \del_in_imag_pl_d~6 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~6 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~6_combout ),
	.cout());
defparam \del_in_real_pl_d~6 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[6]~6 (
	.dataa(out_real_61),
	.datab(out_imag_61),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[6]~6_combout ),
	.cout());
defparam \in_real_cmm[6]~6 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[7]~7 (
	.dataa(out_imag_71),
	.datab(out_real_71),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[7]~7_combout ),
	.cout());
defparam \in_imag_cmm[7]~7 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[7]~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~7 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~7_combout ),
	.cout());
defparam \del_in_imag_pl_d~7 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][7] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~7 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~7_combout ),
	.cout());
defparam \del_in_real_pl_d~7 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[7]~7 (
	.dataa(out_real_71),
	.datab(out_imag_71),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[7]~7_combout ),
	.cout());
defparam \in_real_cmm[7]~7 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_cmm[8]~8 (
	.dataa(out_imag_81),
	.datab(out_real_81),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_imag_cmm[8]~8_combout ),
	.cout());
defparam \in_imag_cmm[8]~8 .lut_mask = 16'hEFFE;
defparam \in_imag_cmm[8]~8 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_cmm_d[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] .power_up = "low";

cycloneiv_lcell_comb \del_in_imag_pl_d~8 (
	.dataa(\generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ),
	.datab(\generate_delay_less_pipeline:in_imag_cmm_d[8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_imag_pl_d~8_combout ),
	.cout());
defparam \del_in_imag_pl_d~8 .lut_mask = 16'hAACC;
defparam \del_in_imag_pl_d~8 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_cmm_d[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][9] .power_up = "low";

cycloneiv_lcell_comb \del_in_real_pl_d~8 (
	.dataa(\generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ),
	.datab(\generate_delay_less_pipeline:in_real_cmm_d[8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\del_in_real_pl_d~8_combout ),
	.cout());
defparam \del_in_real_pl_d~8 .lut_mask = 16'hAACC;
defparam \del_in_real_pl_d~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_cmm[8]~8 (
	.dataa(out_real_81),
	.datab(out_imag_81),
	.datac(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\in_real_cmm[8]~8_combout ),
	.cout());
defparam \in_real_cmm[8]~8 .lut_mask = 16'hEFFE;
defparam \in_real_cmm[8]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb cmm_control(
	.dataa(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\bf_control_inst|bf_counter_inst|control_s[2]~q ),
	.cin(gnd),
	.combout(\cmm_control~combout ),
	.cout());
defparam cmm_control.lut_mask = 16'hAAFF;
defparam cmm_control.sum_lutc_input = "datac";

dffeas \out_imag[2] (
	.clk(clk),
	.d(\out_imag~0_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_2),
	.prn(vcc));
defparam \out_imag[2] .is_wysiwyg = "true";
defparam \out_imag[2] .power_up = "low";

dffeas \out_real[2] (
	.clk(clk),
	.d(\out_real~0_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_2),
	.prn(vcc));
defparam \out_real[2] .is_wysiwyg = "true";
defparam \out_real[2] .power_up = "low";

dffeas \out_imag[3] (
	.clk(clk),
	.d(\out_imag~1_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_3),
	.prn(vcc));
defparam \out_imag[3] .is_wysiwyg = "true";
defparam \out_imag[3] .power_up = "low";

dffeas \out_real[3] (
	.clk(clk),
	.d(\out_real~1_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_3),
	.prn(vcc));
defparam \out_real[3] .is_wysiwyg = "true";
defparam \out_real[3] .power_up = "low";

dffeas \out_imag[4] (
	.clk(clk),
	.d(\out_imag~2_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_4),
	.prn(vcc));
defparam \out_imag[4] .is_wysiwyg = "true";
defparam \out_imag[4] .power_up = "low";

dffeas \out_real[4] (
	.clk(clk),
	.d(\out_real~2_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_4),
	.prn(vcc));
defparam \out_real[4] .is_wysiwyg = "true";
defparam \out_real[4] .power_up = "low";

dffeas \out_imag[5] (
	.clk(clk),
	.d(\out_imag~3_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_5),
	.prn(vcc));
defparam \out_imag[5] .is_wysiwyg = "true";
defparam \out_imag[5] .power_up = "low";

dffeas \out_real[5] (
	.clk(clk),
	.d(\out_real~3_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_5),
	.prn(vcc));
defparam \out_real[5] .is_wysiwyg = "true";
defparam \out_real[5] .power_up = "low";

dffeas \out_imag[6] (
	.clk(clk),
	.d(\out_imag~4_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_6),
	.prn(vcc));
defparam \out_imag[6] .is_wysiwyg = "true";
defparam \out_imag[6] .power_up = "low";

dffeas \out_real[6] (
	.clk(clk),
	.d(\out_real~4_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_6),
	.prn(vcc));
defparam \out_real[6] .is_wysiwyg = "true";
defparam \out_real[6] .power_up = "low";

dffeas \out_imag[7] (
	.clk(clk),
	.d(\out_imag~5_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_7),
	.prn(vcc));
defparam \out_imag[7] .is_wysiwyg = "true";
defparam \out_imag[7] .power_up = "low";

dffeas \out_real[7] (
	.clk(clk),
	.d(\out_real~5_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_7),
	.prn(vcc));
defparam \out_real[7] .is_wysiwyg = "true";
defparam \out_real[7] .power_up = "low";

dffeas \out_imag[8] (
	.clk(clk),
	.d(\out_imag~6_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_8),
	.prn(vcc));
defparam \out_imag[8] .is_wysiwyg = "true";
defparam \out_imag[8] .power_up = "low";

dffeas \out_real[8] (
	.clk(clk),
	.d(\out_real~6_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_8),
	.prn(vcc));
defparam \out_real[8] .is_wysiwyg = "true";
defparam \out_real[8] .power_up = "low";

dffeas \out_imag[9] (
	.clk(clk),
	.d(\out_imag~7_combout ),
	.asdata(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_imag_9),
	.prn(vcc));
defparam \out_imag[9] .is_wysiwyg = "true";
defparam \out_imag[9] .power_up = "low";

dffeas \out_real[9] (
	.clk(clk),
	.d(\out_real~7_combout ),
	.asdata(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(\s_sel_d[1]~q ),
	.ena(enable),
	.q(out_real_9),
	.prn(vcc));
defparam \out_real[9] .is_wysiwyg = "true";
defparam \out_real[9] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\out_valid_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

dffeas out_eop(
	.clk(clk),
	.d(\out_eop_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_eop1),
	.prn(vcc));
defparam out_eop.is_wysiwyg = "true";
defparam out_eop.power_up = "low";

dffeas out_sop(
	.clk(clk),
	.d(\out_sop_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_sop1),
	.prn(vcc));
defparam out_sop.is_wysiwyg = "true";
defparam out_sop.power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][2] .power_up = "low";

cycloneiv_lcell_comb \out_imag~0 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~0_combout ),
	.cout());
defparam \out_imag~0 .lut_mask = 16'hAACC;
defparam \out_imag~0 .sum_lutc_input = "datac";

dffeas \s_sel_d[0] (
	.clk(clk),
	.d(\bf_control_inst|bf_counter_inst|control_s[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[0]~q ),
	.prn(vcc));
defparam \s_sel_d[0] .is_wysiwyg = "true";
defparam \s_sel_d[0] .power_up = "low";

dffeas \s_sel_d[1] (
	.clk(clk),
	.d(\s_sel_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[1]~q ),
	.prn(vcc));
defparam \s_sel_d[1] .is_wysiwyg = "true";
defparam \s_sel_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][2] .power_up = "low";

cycloneiv_lcell_comb \out_real~0 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~0_combout ),
	.cout());
defparam \out_real~0 .lut_mask = 16'hAACC;
defparam \out_real~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][3] .power_up = "low";

cycloneiv_lcell_comb \out_imag~1 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~1_combout ),
	.cout());
defparam \out_imag~1 .lut_mask = 16'hAACC;
defparam \out_imag~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][3] .power_up = "low";

cycloneiv_lcell_comb \out_real~1 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~1_combout ),
	.cout());
defparam \out_real~1 .lut_mask = 16'hAACC;
defparam \out_real~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][4] .power_up = "low";

cycloneiv_lcell_comb \out_imag~2 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~2_combout ),
	.cout());
defparam \out_imag~2 .lut_mask = 16'hAACC;
defparam \out_imag~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][4] .power_up = "low";

cycloneiv_lcell_comb \out_real~2 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~2_combout ),
	.cout());
defparam \out_real~2 .lut_mask = 16'hAACC;
defparam \out_real~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][5] .power_up = "low";

cycloneiv_lcell_comb \out_imag~3 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~3_combout ),
	.cout());
defparam \out_imag~3 .lut_mask = 16'hAACC;
defparam \out_imag~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][5] .power_up = "low";

cycloneiv_lcell_comb \out_real~3 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~3_combout ),
	.cout());
defparam \out_real~3 .lut_mask = 16'hAACC;
defparam \out_real~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][6] .power_up = "low";

cycloneiv_lcell_comb \out_imag~4 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~4_combout ),
	.cout());
defparam \out_imag~4 .lut_mask = 16'hAACC;
defparam \out_imag~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][6] .power_up = "low";

cycloneiv_lcell_comb \out_real~4 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~4_combout ),
	.cout());
defparam \out_real~4 .lut_mask = 16'hAACC;
defparam \out_real~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][7] .power_up = "low";

cycloneiv_lcell_comb \out_imag~5 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~5_combout ),
	.cout());
defparam \out_imag~5 .lut_mask = 16'hAACC;
defparam \out_imag~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][7] .power_up = "low";

cycloneiv_lcell_comb \out_real~5 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~5_combout ),
	.cout());
defparam \out_real~5 .lut_mask = 16'hAACC;
defparam \out_real~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][8] .power_up = "low";

cycloneiv_lcell_comb \out_imag~6 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~6_combout ),
	.cout());
defparam \out_imag~6 .lut_mask = 16'hAACC;
defparam \out_imag~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][8] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][8] .power_up = "low";

cycloneiv_lcell_comb \out_real~6 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~6_combout ),
	.cout());
defparam \out_real~6 .lut_mask = 16'hAACC;
defparam \out_real~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][9] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][9] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[1][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[1][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[1][9] .power_up = "low";

cycloneiv_lcell_comb \out_imag~7 (
	.dataa(\generate_delay_less_pipeline:adder2_out_imag_d[1][9]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_imag~7_combout ),
	.cout());
defparam \out_imag~7 .lut_mask = 16'hAACC;
defparam \out_imag~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][9] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][9] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[1][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[1][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[1][9] .power_up = "low";

cycloneiv_lcell_comb \out_real~7 (
	.dataa(\generate_delay_less_pipeline:adder2_out_real_d[1][9]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ),
	.datac(gnd),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\out_real~7_combout ),
	.cout());
defparam \out_real~7 .lut_mask = 16'hAACC;
defparam \out_real~7 .sum_lutc_input = "datac";

dffeas \out_valid_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_valid~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[0]~q ),
	.prn(vcc));
defparam \out_valid_d[0] .is_wysiwyg = "true";
defparam \out_valid_d[0] .power_up = "low";

dffeas \out_valid_d[1] (
	.clk(clk),
	.d(\out_valid_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[1]~q ),
	.prn(vcc));
defparam \out_valid_d[1] .is_wysiwyg = "true";
defparam \out_valid_d[1] .power_up = "low";

dffeas \out_inverse_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_inverse~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_inverse_d[0]~q ),
	.prn(vcc));
defparam \out_inverse_d[0] .is_wysiwyg = "true";
defparam \out_inverse_d[0] .power_up = "low";

dffeas \out_eop_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_eop~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_eop_d[0]~q ),
	.prn(vcc));
defparam \out_eop_d[0] .is_wysiwyg = "true";
defparam \out_eop_d[0] .power_up = "low";

dffeas \out_sop_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_sop~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_sop_d[0]~q ),
	.prn(vcc));
defparam \out_sop_d[0] .is_wysiwyg = "true";
defparam \out_sop_d[0] .power_up = "low";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_4 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	t_sel_d,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	t_sel_d;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_5 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.t_sel_d(t_sel_d),
	.generate_delay_less_pipelinein_imag_cmm_d2(generate_delay_less_pipelinein_imag_cmm_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.generate_delay_less_pipelinein_imag_cmm_d1(generate_delay_less_pipelinein_imag_cmm_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.generate_delay_less_pipelinein_imag_cmm_d0(generate_delay_less_pipelinein_imag_cmm_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.generate_delay_less_pipelinein_imag_cmm_d3(generate_delay_less_pipelinein_imag_cmm_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.generate_delay_less_pipelinein_imag_cmm_d4(generate_delay_less_pipelinein_imag_cmm_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.generate_delay_less_pipelinein_imag_cmm_d5(generate_delay_less_pipelinein_imag_cmm_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.generate_delay_less_pipelinein_imag_cmm_d6(generate_delay_less_pipelinein_imag_cmm_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.generate_delay_less_pipelinein_imag_cmm_d7(generate_delay_less_pipelinein_imag_cmm_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.generate_delay_less_pipelinein_imag_cmm_d8(generate_delay_less_pipelinein_imag_cmm_d8),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_5 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	t_sel_d,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	t_sel_d;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.t_sel_d(t_sel_d),
	.generate_delay_less_pipelinein_imag_cmm_d2(generate_delay_less_pipelinein_imag_cmm_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.generate_delay_less_pipelinein_imag_cmm_d1(generate_delay_less_pipelinein_imag_cmm_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.generate_delay_less_pipelinein_imag_cmm_d0(generate_delay_less_pipelinein_imag_cmm_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.generate_delay_less_pipelinein_imag_cmm_d3(generate_delay_less_pipelinein_imag_cmm_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.generate_delay_less_pipelinein_imag_cmm_d4(generate_delay_less_pipelinein_imag_cmm_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.generate_delay_less_pipelinein_imag_cmm_d5(generate_delay_less_pipelinein_imag_cmm_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.generate_delay_less_pipelinein_imag_cmm_d6(generate_delay_less_pipelinein_imag_cmm_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.generate_delay_less_pipelinein_imag_cmm_d7(generate_delay_less_pipelinein_imag_cmm_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.generate_delay_less_pipelinein_imag_cmm_d8(generate_delay_less_pipelinein_imag_cmm_d8),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	t_sel_d,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	t_sel_d;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d2),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d1),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d0),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(t_sel_d),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h00BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d3),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d4),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d5),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d6),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d7),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(t_sel_d),
	.datad(generate_delay_less_pipelinein_imag_cmm_d8),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_5 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_6 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d12(generate_delay_less_pipelinedel_in_real_pl_d12),
	.generate_delay_less_pipelinein_real_cmm_d2(generate_delay_less_pipelinein_real_cmm_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d11(generate_delay_less_pipelinedel_in_real_pl_d11),
	.generate_delay_less_pipelinein_real_cmm_d1(generate_delay_less_pipelinein_real_cmm_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d10(generate_delay_less_pipelinedel_in_real_pl_d10),
	.generate_delay_less_pipelinein_real_cmm_d0(generate_delay_less_pipelinein_real_cmm_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d13(generate_delay_less_pipelinedel_in_real_pl_d13),
	.generate_delay_less_pipelinein_real_cmm_d3(generate_delay_less_pipelinein_real_cmm_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d14(generate_delay_less_pipelinedel_in_real_pl_d14),
	.generate_delay_less_pipelinein_real_cmm_d4(generate_delay_less_pipelinein_real_cmm_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d15(generate_delay_less_pipelinedel_in_real_pl_d15),
	.generate_delay_less_pipelinein_real_cmm_d5(generate_delay_less_pipelinein_real_cmm_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d16(generate_delay_less_pipelinedel_in_real_pl_d16),
	.generate_delay_less_pipelinein_real_cmm_d6(generate_delay_less_pipelinein_real_cmm_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d17(generate_delay_less_pipelinedel_in_real_pl_d17),
	.generate_delay_less_pipelinein_real_cmm_d7(generate_delay_less_pipelinein_real_cmm_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d18(generate_delay_less_pipelinedel_in_real_pl_d18),
	.generate_delay_less_pipelinein_real_cmm_d8(generate_delay_less_pipelinein_real_cmm_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_6 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_1 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d12(generate_delay_less_pipelinedel_in_real_pl_d12),
	.generate_delay_less_pipelinein_real_cmm_d2(generate_delay_less_pipelinein_real_cmm_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d11(generate_delay_less_pipelinedel_in_real_pl_d11),
	.generate_delay_less_pipelinein_real_cmm_d1(generate_delay_less_pipelinein_real_cmm_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d10(generate_delay_less_pipelinedel_in_real_pl_d10),
	.generate_delay_less_pipelinein_real_cmm_d0(generate_delay_less_pipelinein_real_cmm_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d13(generate_delay_less_pipelinedel_in_real_pl_d13),
	.generate_delay_less_pipelinein_real_cmm_d3(generate_delay_less_pipelinein_real_cmm_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d14(generate_delay_less_pipelinedel_in_real_pl_d14),
	.generate_delay_less_pipelinein_real_cmm_d4(generate_delay_less_pipelinein_real_cmm_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d15(generate_delay_less_pipelinedel_in_real_pl_d15),
	.generate_delay_less_pipelinein_real_cmm_d5(generate_delay_less_pipelinein_real_cmm_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d16(generate_delay_less_pipelinedel_in_real_pl_d16),
	.generate_delay_less_pipelinein_real_cmm_d6(generate_delay_less_pipelinein_real_cmm_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d17(generate_delay_less_pipelinedel_in_real_pl_d17),
	.generate_delay_less_pipelinein_real_cmm_d7(generate_delay_less_pipelinein_real_cmm_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d18(generate_delay_less_pipelinedel_in_real_pl_d18),
	.generate_delay_less_pipelinein_real_cmm_d8(generate_delay_less_pipelinein_real_cmm_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_1 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d10),
	.datab(generate_delay_less_pipelinein_real_cmm_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00EE;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d11),
	.datab(generate_delay_less_pipelinein_real_cmm_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h007F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d12),
	.datab(generate_delay_less_pipelinein_real_cmm_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d13),
	.datab(generate_delay_less_pipelinein_real_cmm_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d14),
	.datab(generate_delay_less_pipelinein_real_cmm_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d15),
	.datab(generate_delay_less_pipelinein_real_cmm_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d16),
	.datab(generate_delay_less_pipelinein_real_cmm_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d17),
	.datab(generate_delay_less_pipelinein_real_cmm_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d18),
	.datab(generate_delay_less_pipelinein_real_cmm_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d18),
	.datab(generate_delay_less_pipelinein_real_cmm_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_6 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	cmm_control_d,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	cmm_control_d;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_7 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinein_imag_cmm_d2(generate_delay_less_pipelinein_imag_cmm_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.generate_delay_less_pipelinein_imag_cmm_d1(generate_delay_less_pipelinein_imag_cmm_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.generate_delay_less_pipelinein_imag_cmm_d0(generate_delay_less_pipelinein_imag_cmm_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.generate_delay_less_pipelinein_imag_cmm_d3(generate_delay_less_pipelinein_imag_cmm_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.generate_delay_less_pipelinein_imag_cmm_d4(generate_delay_less_pipelinein_imag_cmm_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.generate_delay_less_pipelinein_imag_cmm_d5(generate_delay_less_pipelinein_imag_cmm_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.generate_delay_less_pipelinein_imag_cmm_d6(generate_delay_less_pipelinein_imag_cmm_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.generate_delay_less_pipelinein_imag_cmm_d7(generate_delay_less_pipelinein_imag_cmm_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.generate_delay_less_pipelinein_imag_cmm_d8(generate_delay_less_pipelinein_imag_cmm_d8),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.cmm_control_d(cmm_control_d),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_7 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	cmm_control_d,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	cmm_control_d;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_2 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinein_imag_cmm_d2(generate_delay_less_pipelinein_imag_cmm_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d12(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.generate_delay_less_pipelinein_imag_cmm_d1(generate_delay_less_pipelinein_imag_cmm_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d11(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.generate_delay_less_pipelinein_imag_cmm_d0(generate_delay_less_pipelinein_imag_cmm_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d10(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.generate_delay_less_pipelinein_imag_cmm_d3(generate_delay_less_pipelinein_imag_cmm_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d13(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.generate_delay_less_pipelinein_imag_cmm_d4(generate_delay_less_pipelinein_imag_cmm_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d14(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.generate_delay_less_pipelinein_imag_cmm_d5(generate_delay_less_pipelinein_imag_cmm_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d15(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.generate_delay_less_pipelinein_imag_cmm_d6(generate_delay_less_pipelinein_imag_cmm_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d16(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.generate_delay_less_pipelinein_imag_cmm_d7(generate_delay_less_pipelinein_imag_cmm_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d17(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.generate_delay_less_pipelinein_imag_cmm_d8(generate_delay_less_pipelinein_imag_cmm_d8),
	.generate_delay_less_pipelinedel_in_imag_pl_d18(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.cmm_control_d(cmm_control_d),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_2 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinein_imag_cmm_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d12,
	generate_delay_less_pipelinein_imag_cmm_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d11,
	generate_delay_less_pipelinein_imag_cmm_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d10,
	generate_delay_less_pipelinein_imag_cmm_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d13,
	generate_delay_less_pipelinein_imag_cmm_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d14,
	generate_delay_less_pipelinein_imag_cmm_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d15,
	generate_delay_less_pipelinein_imag_cmm_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d16,
	generate_delay_less_pipelinein_imag_cmm_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d17,
	generate_delay_less_pipelinein_imag_cmm_d8,
	generate_delay_less_pipelinedel_in_imag_pl_d18,
	cmm_control_d,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinein_imag_cmm_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d12;
input 	generate_delay_less_pipelinein_imag_cmm_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d11;
input 	generate_delay_less_pipelinein_imag_cmm_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d10;
input 	generate_delay_less_pipelinein_imag_cmm_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d13;
input 	generate_delay_less_pipelinein_imag_cmm_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d14;
input 	generate_delay_less_pipelinein_imag_cmm_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d15;
input 	generate_delay_less_pipelinein_imag_cmm_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d16;
input 	generate_delay_less_pipelinein_imag_cmm_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d17;
input 	generate_delay_less_pipelinein_imag_cmm_d8;
input 	generate_delay_less_pipelinedel_in_imag_pl_d18;
input 	cmm_control_d;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d2),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d1),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d0),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(cmm_control_d),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h0055;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~2_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d10),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h00BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~1_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d11),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .lut_mask = 16'h00DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~0_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d12),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d3),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~3_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d13),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d4),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~4_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d14),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d5),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~5_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d15),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d6),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~6_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d16),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d7),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~7_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d17),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(generate_delay_less_pipelinein_imag_cmm_d8),
	.datad(cmm_control_d),
	.cin(gnd),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 .lut_mask = 16'h0FF0;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~26 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 (
	.dataa(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|_~8_combout ),
	.datab(generate_delay_less_pipelinedel_in_imag_pl_d18),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~27 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~28 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_7 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_8 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d12(generate_delay_less_pipelinedel_in_real_pl_d12),
	.generate_delay_less_pipelinein_real_cmm_d2(generate_delay_less_pipelinein_real_cmm_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d11(generate_delay_less_pipelinedel_in_real_pl_d11),
	.generate_delay_less_pipelinein_real_cmm_d1(generate_delay_less_pipelinein_real_cmm_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d10(generate_delay_less_pipelinedel_in_real_pl_d10),
	.generate_delay_less_pipelinein_real_cmm_d0(generate_delay_less_pipelinein_real_cmm_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d13(generate_delay_less_pipelinedel_in_real_pl_d13),
	.generate_delay_less_pipelinein_real_cmm_d3(generate_delay_less_pipelinein_real_cmm_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d14(generate_delay_less_pipelinedel_in_real_pl_d14),
	.generate_delay_less_pipelinein_real_cmm_d4(generate_delay_less_pipelinein_real_cmm_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d15(generate_delay_less_pipelinedel_in_real_pl_d15),
	.generate_delay_less_pipelinein_real_cmm_d5(generate_delay_less_pipelinein_real_cmm_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d16(generate_delay_less_pipelinedel_in_real_pl_d16),
	.generate_delay_less_pipelinein_real_cmm_d6(generate_delay_less_pipelinein_real_cmm_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d17(generate_delay_less_pipelinedel_in_real_pl_d17),
	.generate_delay_less_pipelinein_real_cmm_d7(generate_delay_less_pipelinein_real_cmm_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d18(generate_delay_less_pipelinedel_in_real_pl_d18),
	.generate_delay_less_pipelinein_real_cmm_d8(generate_delay_less_pipelinein_real_cmm_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_8 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_3 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d12(generate_delay_less_pipelinedel_in_real_pl_d12),
	.generate_delay_less_pipelinein_real_cmm_d2(generate_delay_less_pipelinein_real_cmm_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d11(generate_delay_less_pipelinedel_in_real_pl_d11),
	.generate_delay_less_pipelinein_real_cmm_d1(generate_delay_less_pipelinein_real_cmm_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d10(generate_delay_less_pipelinedel_in_real_pl_d10),
	.generate_delay_less_pipelinein_real_cmm_d0(generate_delay_less_pipelinein_real_cmm_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d13(generate_delay_less_pipelinedel_in_real_pl_d13),
	.generate_delay_less_pipelinein_real_cmm_d3(generate_delay_less_pipelinein_real_cmm_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d14(generate_delay_less_pipelinedel_in_real_pl_d14),
	.generate_delay_less_pipelinein_real_cmm_d4(generate_delay_less_pipelinein_real_cmm_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d15(generate_delay_less_pipelinedel_in_real_pl_d15),
	.generate_delay_less_pipelinein_real_cmm_d5(generate_delay_less_pipelinein_real_cmm_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d16(generate_delay_less_pipelinedel_in_real_pl_d16),
	.generate_delay_less_pipelinein_real_cmm_d6(generate_delay_less_pipelinein_real_cmm_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d17(generate_delay_less_pipelinedel_in_real_pl_d17),
	.generate_delay_less_pipelinein_real_cmm_d7(generate_delay_less_pipelinein_real_cmm_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d18(generate_delay_less_pipelinedel_in_real_pl_d18),
	.generate_delay_less_pipelinein_real_cmm_d8(generate_delay_less_pipelinein_real_cmm_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_3 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d12,
	generate_delay_less_pipelinein_real_cmm_d2,
	generate_delay_less_pipelinedel_in_real_pl_d11,
	generate_delay_less_pipelinein_real_cmm_d1,
	generate_delay_less_pipelinedel_in_real_pl_d10,
	generate_delay_less_pipelinein_real_cmm_d0,
	generate_delay_less_pipelinedel_in_real_pl_d13,
	generate_delay_less_pipelinein_real_cmm_d3,
	generate_delay_less_pipelinedel_in_real_pl_d14,
	generate_delay_less_pipelinein_real_cmm_d4,
	generate_delay_less_pipelinedel_in_real_pl_d15,
	generate_delay_less_pipelinein_real_cmm_d5,
	generate_delay_less_pipelinedel_in_real_pl_d16,
	generate_delay_less_pipelinein_real_cmm_d6,
	generate_delay_less_pipelinedel_in_real_pl_d17,
	generate_delay_less_pipelinein_real_cmm_d7,
	generate_delay_less_pipelinedel_in_real_pl_d18,
	generate_delay_less_pipelinein_real_cmm_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d12;
input 	generate_delay_less_pipelinein_real_cmm_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d11;
input 	generate_delay_less_pipelinein_real_cmm_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d10;
input 	generate_delay_less_pipelinein_real_cmm_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d13;
input 	generate_delay_less_pipelinein_real_cmm_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d14;
input 	generate_delay_less_pipelinein_real_cmm_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d15;
input 	generate_delay_less_pipelinein_real_cmm_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d16;
input 	generate_delay_less_pipelinein_real_cmm_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d17;
input 	generate_delay_less_pipelinein_real_cmm_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d18;
input 	generate_delay_less_pipelinein_real_cmm_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d10),
	.datab(generate_delay_less_pipelinein_real_cmm_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00BB;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d11),
	.datab(generate_delay_less_pipelinein_real_cmm_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h00DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d12),
	.datab(generate_delay_less_pipelinein_real_cmm_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d13),
	.datab(generate_delay_less_pipelinein_real_cmm_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d14),
	.datab(generate_delay_less_pipelinein_real_cmm_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d15),
	.datab(generate_delay_less_pipelinein_real_cmm_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d16),
	.datab(generate_delay_less_pipelinein_real_cmm_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d17),
	.datab(generate_delay_less_pipelinein_real_cmm_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d18),
	.datab(generate_delay_less_pipelinein_real_cmm_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d18),
	.datab(generate_delay_less_pipelinein_real_cmm_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:0:r22_stage|gen_bfii:bfii_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_bf_control_1 (
	out_control_2,
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	control_s_1,
	out_valid1,
	out_inverse1,
	out_eop1,
	out_sop1,
	out_valid2,
	control_s_2,
	out_inverse2,
	out_sop2,
	out_control_1,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	out_control_2;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
input 	fftpts_less_one_0;
input 	fftpts_less_one_1;
input 	fftpts_less_one_2;
input 	fftpts_less_one_3;
output 	control_s_1;
output 	out_valid1;
output 	out_inverse1;
output 	out_eop1;
input 	out_sop1;
input 	out_valid2;
output 	control_s_2;
input 	out_inverse2;
output 	out_sop2;
output 	out_control_1;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \bf_counter_inst|counter_p~0_combout ;
wire \Add0~0_combout ;
wire \Equal0~0_combout ;
wire \Add3~1_combout ;
wire \in_cnt~3_combout ;
wire \in_cnt[2]~q ;
wire \Add3~0_combout ;
wire \in_cnt~2_combout ;
wire \in_cnt[3]~q ;
wire \Equal0~1_combout ;
wire \in_cnt~1_combout ;
wire \in_cnt[0]~q ;
wire \in_cnt~0_combout ;
wire \in_cnt[1]~q ;
wire \Equal1~0_combout ;
wire \Add4~1_combout ;
wire \out_cnt[2]~5_combout ;
wire \out_cnt[2]~q ;
wire \Add4~0_combout ;
wire \out_cnt[3]~4_combout ;
wire \out_cnt[3]~q ;
wire \Equal2~1_combout ;
wire \out_eop~0_combout ;
wire \out_cnt[0]~3_combout ;
wire \out_cnt[0]~q ;
wire \out_cnt[0]~0_combout ;
wire \Equal1~1_combout ;
wire \out_cnt[3]~1_combout ;
wire \out_cnt[1]~2_combout ;
wire \out_cnt[1]~q ;
wire \Equal2~0_combout ;
wire \Equal2~2_combout ;
wire \shift~4_combout ;
wire \shift~q ;
wire \out_inverse~0_combout ;


ifft_8p_auk_dspip_r22sdf_counter_1 bf_counter_inst(
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.control_s_1(control_s_1),
	.out_sop(out_sop1),
	.out_valid(out_valid2),
	.counter_p(\bf_counter_inst|counter_p~0_combout ),
	.control_s_2(control_s_2),
	.out_control_1(out_control_1),
	.clk(clk),
	.reset(reset));

dffeas \out_control[2] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(out_control_1),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(curr_pwr_2_s),
	.ena(enable),
	.q(out_control_2),
	.prn(vcc));
defparam \out_control[2] .is_wysiwyg = "true";
defparam \out_control[2] .power_up = "low";

cycloneiv_lcell_comb out_valid(
	.dataa(\shift~q ),
	.datab(control_s_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'hEEEE;
defparam out_valid.sum_lutc_input = "datac";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

dffeas out_eop(
	.clk(clk),
	.d(\out_eop~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_eop1),
	.prn(vcc));
defparam out_eop.is_wysiwyg = "true";
defparam out_eop.power_up = "low";

dffeas out_sop(
	.clk(clk),
	.d(\Equal1~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_sop2),
	.prn(vcc));
defparam out_sop.is_wysiwyg = "true";
defparam out_sop.power_up = "low";

dffeas \out_control[1] (
	.clk(clk),
	.d(vcc),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_control_1),
	.prn(vcc));
defparam \out_control[1] .is_wysiwyg = "true";
defparam \out_control[1] .power_up = "low";

cycloneiv_lcell_comb \Add0~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(curr_pwr_2_s),
	.datad(out_control_1),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
defparam \Add0~0 .lut_mask = 16'h0FF0;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\in_cnt[1]~q ),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(\in_cnt[2]~q ),
	.datac(\in_cnt[0]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'hC33C;
defparam \Add3~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~3 (
	.dataa(\Add3~1_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~3_combout ),
	.cout());
defparam \in_cnt~3 .lut_mask = 16'hAFFF;
defparam \in_cnt~3 .sum_lutc_input = "datac";

dffeas \in_cnt[2] (
	.clk(clk),
	.d(\in_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[2]~q ),
	.prn(vcc));
defparam \in_cnt[2] .is_wysiwyg = "true";
defparam \in_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Add3~0 (
	.dataa(\in_cnt[3]~q ),
	.datab(\in_cnt[2]~q ),
	.datac(\in_cnt[0]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h6996;
defparam \Add3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~2 (
	.dataa(\Add3~0_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~2_combout ),
	.cout());
defparam \in_cnt~2 .lut_mask = 16'hAFFF;
defparam \in_cnt~2 .sum_lutc_input = "datac";

dffeas \in_cnt[3] (
	.clk(clk),
	.d(\in_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[3]~q ),
	.prn(vcc));
defparam \in_cnt[3] .is_wysiwyg = "true";
defparam \in_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \Equal0~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\in_cnt[3]~q ),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~1 (
	.dataa(\in_cnt[0]~q ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_cnt~1_combout ),
	.cout());
defparam \in_cnt~1 .lut_mask = 16'h7F7F;
defparam \in_cnt~1 .sum_lutc_input = "datac";

dffeas \in_cnt[0] (
	.clk(clk),
	.d(\in_cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[0]~q ),
	.prn(vcc));
defparam \in_cnt[0] .is_wysiwyg = "true";
defparam \in_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \in_cnt~0 (
	.dataa(\in_cnt[0]~q ),
	.datab(\in_cnt[1]~q ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~0_combout ),
	.cout());
defparam \in_cnt~0 .lut_mask = 16'h6FFF;
defparam \in_cnt~0 .sum_lutc_input = "datac";

dffeas \in_cnt[1] (
	.clk(clk),
	.d(\in_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[1]~q ),
	.prn(vcc));
defparam \in_cnt[1] .is_wysiwyg = "true";
defparam \in_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal1~0 (
	.dataa(curr_pwr_2_s),
	.datab(\in_cnt[1]~q ),
	.datac(\in_cnt[0]~q ),
	.datad(\in_cnt[3]~q ),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'h96FF;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(\out_cnt[2]~q ),
	.datac(\out_cnt[0]~q ),
	.datad(\out_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add4~1_combout ),
	.cout());
defparam \Add4~1 .lut_mask = 16'hC33C;
defparam \Add4~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[2]~5 (
	.dataa(\out_cnt[2]~q ),
	.datab(\out_cnt[3]~1_combout ),
	.datac(\Add4~1_combout ),
	.datad(\out_eop~0_combout ),
	.cin(gnd),
	.combout(\out_cnt[2]~5_combout ),
	.cout());
defparam \out_cnt[2]~5 .lut_mask = 16'hB8FF;
defparam \out_cnt[2]~5 .sum_lutc_input = "datac";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Add4~0 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[0]~q ),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout());
defparam \Add4~0 .lut_mask = 16'h6996;
defparam \Add4~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~4 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[3]~1_combout ),
	.datac(\Add4~0_combout ),
	.datad(\out_eop~0_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~4_combout ),
	.cout());
defparam \out_cnt[3]~4 .lut_mask = 16'hB8FF;
defparam \out_cnt[3]~4 .sum_lutc_input = "datac";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \Equal2~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\out_cnt[3]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'h6996;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_eop~0 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\in_cnt[2]~q ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\out_eop~0_combout ),
	.cout());
defparam \out_eop~0 .lut_mask = 16'hFEFF;
defparam \out_eop~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[0]~3 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[3]~1_combout ),
	.datac(gnd),
	.datad(\out_eop~0_combout ),
	.cin(gnd),
	.combout(\out_cnt[0]~3_combout ),
	.cout());
defparam \out_cnt[0]~3 .lut_mask = 16'h66FF;
defparam \out_cnt[0]~3 .sum_lutc_input = "datac";

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \out_cnt[0]~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\out_cnt[0]~0_combout ),
	.cout());
defparam \out_cnt[0]~0 .lut_mask = 16'h7FFF;
defparam \out_cnt[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal1~1 (
	.dataa(\Equal1~0_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
defparam \Equal1~1 .lut_mask = 16'hAAFF;
defparam \Equal1~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~1 (
	.dataa(enable),
	.datab(\out_cnt[0]~0_combout ),
	.datac(\Equal2~2_combout ),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~1_combout ),
	.cout());
defparam \out_cnt[3]~1 .lut_mask = 16'hDFFF;
defparam \out_cnt[3]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[1]~2 (
	.dataa(\out_cnt[1]~q ),
	.datab(\out_cnt[3]~1_combout ),
	.datac(\out_cnt[0]~q ),
	.datad(\out_eop~0_combout ),
	.cin(gnd),
	.combout(\out_cnt[1]~2_combout ),
	.cout());
defparam \out_cnt[1]~2 .lut_mask = 16'h96FF;
defparam \out_cnt[1]~2 .sum_lutc_input = "datac";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal2~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h6996;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Equal2~2 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
defparam \Equal2~2 .lut_mask = 16'hEEEE;
defparam \Equal2~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shift~4 (
	.dataa(\Equal1~0_combout ),
	.datab(\in_cnt[2]~q ),
	.datac(\shift~q ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(\shift~4_combout ),
	.cout());
defparam \shift~4 .lut_mask = 16'hFBFF;
defparam \shift~4 .sum_lutc_input = "datac";

dffeas shift(
	.clk(clk),
	.d(\shift~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\shift~q ),
	.prn(vcc));
defparam shift.is_wysiwyg = "true";
defparam shift.power_up = "low";

cycloneiv_lcell_comb \out_inverse~0 (
	.dataa(out_inverse1),
	.datab(out_inverse2),
	.datac(\Equal1~1_combout ),
	.datad(enable),
	.cin(gnd),
	.combout(\out_inverse~0_combout ),
	.cout());
defparam \out_inverse~0 .lut_mask = 16'hEFFE;
defparam \out_inverse~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_counter_1 (
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	control_s_1,
	out_sop,
	out_valid,
	counter_p,
	control_s_2,
	out_control_1,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
output 	control_s_1;
input 	out_sop;
input 	out_valid;
output 	counter_p;
output 	control_s_2;
input 	out_control_1;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_s~1_combout ;
wire \control_s[0]~q ;
wire \control_s~0_combout ;
wire \control_s~2_combout ;
wire \control_s~3_combout ;


dffeas \control_s[1] (
	.clk(clk),
	.d(\control_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(counter_p),
	.q(control_s_1),
	.prn(vcc));
defparam \control_s[1] .is_wysiwyg = "true";
defparam \control_s[1] .power_up = "low";

cycloneiv_lcell_comb \counter_p~0 (
	.dataa(out_valid),
	.datab(out_valid_s),
	.datac(sop),
	.datad(out_stall_d),
	.cin(gnd),
	.combout(counter_p),
	.cout());
defparam \counter_p~0 .lut_mask = 16'hACFF;
defparam \counter_p~0 .sum_lutc_input = "datac";

dffeas \control_s[2] (
	.clk(clk),
	.d(\control_s~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(counter_p),
	.q(control_s_2),
	.prn(vcc));
defparam \control_s[2] .is_wysiwyg = "true";
defparam \control_s[2] .power_up = "low";

cycloneiv_lcell_comb \control_s~1 (
	.dataa(curr_pwr_2_s),
	.datab(out_sop),
	.datac(gnd),
	.datad(\control_s[0]~q ),
	.cin(gnd),
	.combout(\control_s~1_combout ),
	.cout());
defparam \control_s~1 .lut_mask = 16'h9966;
defparam \control_s~1 .sum_lutc_input = "datac";

dffeas \control_s[0] (
	.clk(clk),
	.d(\control_s~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(counter_p),
	.q(\control_s[0]~q ),
	.prn(vcc));
defparam \control_s[0] .is_wysiwyg = "true";
defparam \control_s[0] .power_up = "low";

cycloneiv_lcell_comb \control_s~0 (
	.dataa(\control_s[0]~q ),
	.datab(control_s_1),
	.datac(out_sop),
	.datad(curr_pwr_2_s),
	.cin(gnd),
	.combout(\control_s~0_combout ),
	.cout());
defparam \control_s~0 .lut_mask = 16'h6996;
defparam \control_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~2 (
	.dataa(curr_pwr_2_s),
	.datab(\control_s[0]~q ),
	.datac(control_s_2),
	.datad(control_s_1),
	.cin(gnd),
	.combout(\control_s~2_combout ),
	.cout());
defparam \control_s~2 .lut_mask = 16'h6996;
defparam \control_s~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~3 (
	.dataa(out_control_1),
	.datab(\control_s~2_combout ),
	.datac(gnd),
	.datad(out_sop),
	.cin(gnd),
	.combout(\control_s~3_combout ),
	.cout());
defparam \control_s~3 .lut_mask = 16'hAACC;
defparam \control_s~3 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_stage_1 (
	stg_imag_next_0,
	stg_real_next_0,
	stg_imag_next_1,
	stg_real_next_1,
	stg_imag_next_2,
	stg_real_next_2,
	stg_imag_next_3,
	stg_real_next_3,
	stg_imag_next_4,
	stg_real_next_4,
	stg_imag_next_5,
	stg_real_next_5,
	stg_imag_next_6,
	stg_real_next_6,
	stg_imag_next_7,
	stg_real_next_7,
	imagtwid_0,
	imagtwid_1,
	imagtwid_2,
	imagtwid_3,
	imagtwid_4,
	imagtwid_5,
	imagtwid_6,
	imagtwid_7,
	curr_blk_s_1,
	out_stall_d,
	out_valid,
	stg_valid_next,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	out_enable,
	processing1,
	out_imag_2,
	out_real_2,
	out_inverse,
	stg_inverse_next,
	out_imag_3,
	out_real_3,
	out_imag_4,
	out_real_4,
	out_imag_5,
	out_real_5,
	out_imag_6,
	out_real_6,
	out_imag_7,
	out_real_7,
	out_imag_8,
	out_real_8,
	out_imag_9,
	out_real_9,
	stg_sop_next,
	stg_eop_next,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	realtwid_0,
	realtwid_1,
	realtwid_2,
	realtwid_3,
	realtwid_4,
	realtwid_5,
	realtwid_6,
	realtwid_7,
	control_s_1,
	control_s_2,
	control_s_0,
	stg_control_next_1,
	stg_control_next_2,
	twid_rd_en,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	stg_imag_next_0;
input 	stg_real_next_0;
input 	stg_imag_next_1;
input 	stg_real_next_1;
input 	stg_imag_next_2;
input 	stg_real_next_2;
input 	stg_imag_next_3;
input 	stg_real_next_3;
input 	stg_imag_next_4;
input 	stg_real_next_4;
input 	stg_imag_next_5;
input 	stg_real_next_5;
input 	stg_imag_next_6;
input 	stg_real_next_6;
input 	stg_imag_next_7;
input 	stg_real_next_7;
input 	imagtwid_0;
input 	imagtwid_1;
input 	imagtwid_2;
input 	imagtwid_3;
input 	imagtwid_4;
input 	imagtwid_5;
input 	imagtwid_6;
input 	imagtwid_7;
input 	curr_blk_s_1;
input 	out_stall_d;
output 	out_valid;
input 	stg_valid_next;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	out_enable;
output 	processing1;
output 	out_imag_2;
output 	out_real_2;
output 	out_inverse;
input 	stg_inverse_next;
output 	out_imag_3;
output 	out_real_3;
output 	out_imag_4;
output 	out_real_4;
output 	out_imag_5;
output 	out_real_5;
output 	out_imag_6;
output 	out_real_6;
output 	out_imag_7;
output 	out_real_7;
output 	out_imag_8;
output 	out_real_8;
output 	out_imag_9;
output 	out_real_9;
input 	stg_sop_next;
input 	stg_eop_next;
input 	fftpts_less_one_0;
input 	fftpts_less_one_1;
input 	fftpts_less_one_2;
input 	fftpts_less_one_3;
input 	realtwid_0;
input 	realtwid_1;
input 	realtwid_2;
input 	realtwid_3;
input 	realtwid_4;
input 	realtwid_5;
input 	realtwid_6;
input 	realtwid_7;
output 	control_s_1;
output 	control_s_2;
output 	control_s_0;
input 	stg_control_next_1;
input 	stg_control_next_2;
output 	twid_rd_en;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[2]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[1]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[0]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[2]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[1]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[0]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[3]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[3]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[4]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[4]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[5]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[5]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[6]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[6]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[7]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[7]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[8]~q ;
wire \gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[8]~q ;
wire \gen_bfi:gen_bfi_only:bfi_inst|out_eop~q ;
wire \gen_cma:cma_inst|out_sop_d[8]~q ;
wire \gen_cma:cma_inst|out_valid_d[8]~q ;
wire \gen_cma:cma_inst|out_inverse_d[8]~q ;
wire \processing_cnt[0]~5_combout ;
wire \processing_cnt[2]~0_combout ;
wire \processing_cnt[2]~1_combout ;
wire \processing_cnt[2]~2_combout ;
wire \processing_cnt[0]~q ;
wire \Add2~2_combout ;
wire \processing_cnt[1]~q ;
wire \Add2~0_combout ;
wire \Add2~1_combout ;
wire \processing_cnt[2]~q ;
wire \res~0_combout ;


ifft_8p_auk_dspip_r22sdf_bfi_1 \gen_bfi:gen_bfi_only:bfi_inst (
	.in_imag({\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[8]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[7]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[6]~q ,
\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[5]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[4]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[3]~q ,
\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[2]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[1]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[0]~q }),
	.in_real({\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[8]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[7]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[6]~q ,
\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[5]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[4]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[3]~q ,
\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[2]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[1]~q ,\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[0]~q }),
	.out_stall_d(out_stall_d),
	.out_valid1(out_valid),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(out_enable),
	.out_imag_2(out_imag_2),
	.out_real_2(out_real_2),
	.out_inverse1(out_inverse),
	.out_imag_3(out_imag_3),
	.out_real_3(out_real_3),
	.out_imag_4(out_imag_4),
	.out_real_4(out_real_4),
	.out_imag_5(out_imag_5),
	.out_real_5(out_real_5),
	.out_imag_6(out_imag_6),
	.out_real_6(out_real_6),
	.out_imag_7(out_imag_7),
	.out_real_7(out_real_7),
	.out_imag_8(out_imag_8),
	.out_real_8(out_real_8),
	.out_imag_9(out_imag_9),
	.out_real_9(out_real_9),
	.out_eop1(\gen_bfi:gen_bfi_only:bfi_inst|out_eop~q ),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.out_sop_d_8(\gen_cma:cma_inst|out_sop_d[8]~q ),
	.out_valid_d_8(\gen_cma:cma_inst|out_valid_d[8]~q ),
	.out_inverse_d_8(\gen_cma:cma_inst|out_inverse_d[8]~q ),
	.clk(clk),
	.reset(reset));

ifft_8p_auk_dspip_r22sdf_cma \gen_cma:cma_inst (
	.stg_imag_next_0(stg_imag_next_0),
	.stg_real_next_0(stg_real_next_0),
	.stg_imag_next_1(stg_imag_next_1),
	.stg_real_next_1(stg_real_next_1),
	.stg_imag_next_2(stg_imag_next_2),
	.stg_real_next_2(stg_real_next_2),
	.stg_imag_next_3(stg_imag_next_3),
	.stg_real_next_3(stg_real_next_3),
	.stg_imag_next_4(stg_imag_next_4),
	.stg_real_next_4(stg_real_next_4),
	.stg_imag_next_5(stg_imag_next_5),
	.stg_real_next_5(stg_real_next_5),
	.stg_imag_next_6(stg_imag_next_6),
	.stg_real_next_6(stg_real_next_6),
	.stg_imag_next_7(stg_imag_next_7),
	.stg_real_next_7(stg_real_next_7),
	.dataout_2(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[2]~q ),
	.dataout_1(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[1]~q ),
	.dataout_0(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[0]~q ),
	.dataout_21(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[2]~q ),
	.dataout_11(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[1]~q ),
	.dataout_01(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[0]~q ),
	.dataout_3(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[3]~q ),
	.dataout_31(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[3]~q ),
	.dataout_4(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[4]~q ),
	.dataout_41(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[4]~q ),
	.dataout_5(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[5]~q ),
	.dataout_51(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[5]~q ),
	.dataout_6(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[6]~q ),
	.dataout_61(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[6]~q ),
	.dataout_7(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[7]~q ),
	.dataout_71(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[7]~q ),
	.dataout_8(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_imag|dataout[8]~q ),
	.dataout_81(\gen_cma:cma_inst|NONA10_C_Mult_Archs:gen_small_mult:round_real|dataout[8]~q ),
	.imagtwid_0(imagtwid_0),
	.imagtwid_1(imagtwid_1),
	.imagtwid_2(imagtwid_2),
	.imagtwid_3(imagtwid_3),
	.imagtwid_4(imagtwid_4),
	.imagtwid_5(imagtwid_5),
	.imagtwid_6(imagtwid_6),
	.imagtwid_7(imagtwid_7),
	.out_stall_d(out_stall_d),
	.stg_valid_next(stg_valid_next),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.out_enable(out_enable),
	.stg_inverse_next(stg_inverse_next),
	.stg_sop_next(stg_sop_next),
	.out_sop_d_8(\gen_cma:cma_inst|out_sop_d[8]~q ),
	.out_valid_d_8(\gen_cma:cma_inst|out_valid_d[8]~q ),
	.out_inverse_d_8(\gen_cma:cma_inst|out_inverse_d[8]~q ),
	.realtwid_0(realtwid_0),
	.realtwid_1(realtwid_1),
	.realtwid_2(realtwid_2),
	.realtwid_3(realtwid_3),
	.realtwid_4(realtwid_4),
	.realtwid_5(realtwid_5),
	.realtwid_6(realtwid_6),
	.realtwid_7(realtwid_7),
	.control_s_1(control_s_1),
	.control_s_2(control_s_2),
	.control_s_0(control_s_0),
	.stg_control_next_1(stg_control_next_1),
	.stg_control_next_2(stg_control_next_2),
	.clk(clk),
	.reset(reset));

dffeas processing(
	.clk(clk),
	.d(\res~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(processing1),
	.prn(vcc));
defparam processing.is_wysiwyg = "true";
defparam processing.power_up = "low";

cycloneiv_lcell_comb \twid_rd_en~0 (
	.dataa(curr_pwr_2_s),
	.datab(stg_valid_next),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(twid_rd_en),
	.cout());
defparam \twid_rd_en~0 .lut_mask = 16'hEEFF;
defparam \twid_rd_en~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[0]~5 (
	.dataa(\processing_cnt[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\processing_cnt[0]~5_combout ),
	.cout());
defparam \processing_cnt[0]~5 .lut_mask = 16'h5555;
defparam \processing_cnt[0]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[2]~0 (
	.dataa(stg_eop_next),
	.datab(curr_pwr_2_s),
	.datac(out_valid),
	.datad(\gen_bfi:gen_bfi_only:bfi_inst|out_eop~q ),
	.cin(gnd),
	.combout(\processing_cnt[2]~0_combout ),
	.cout());
defparam \processing_cnt[2]~0 .lut_mask = 16'h47FF;
defparam \processing_cnt[2]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[2]~1 (
	.dataa(stg_valid_next),
	.datab(stg_sop_next),
	.datac(curr_pwr_2_s),
	.datad(gnd),
	.cin(gnd),
	.combout(\processing_cnt[2]~1_combout ),
	.cout());
defparam \processing_cnt[2]~1 .lut_mask = 16'hB1B1;
defparam \processing_cnt[2]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \processing_cnt[2]~2 (
	.dataa(stg_valid_next),
	.datab(out_enable),
	.datac(\processing_cnt[2]~0_combout ),
	.datad(\processing_cnt[2]~1_combout ),
	.cin(gnd),
	.combout(\processing_cnt[2]~2_combout ),
	.cout());
defparam \processing_cnt[2]~2 .lut_mask = 16'hEFFE;
defparam \processing_cnt[2]~2 .sum_lutc_input = "datac";

dffeas \processing_cnt[0] (
	.clk(clk),
	.d(\processing_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~2_combout ),
	.q(\processing_cnt[0]~q ),
	.prn(vcc));
defparam \processing_cnt[0] .is_wysiwyg = "true";
defparam \processing_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \Add2~2 (
	.dataa(stg_valid_next),
	.datab(stg_sop_next),
	.datac(\processing_cnt[1]~q ),
	.datad(\processing_cnt[0]~q ),
	.cin(gnd),
	.combout(\Add2~2_combout ),
	.cout());
defparam \Add2~2 .lut_mask = 16'h6996;
defparam \Add2~2 .sum_lutc_input = "datac";

dffeas \processing_cnt[1] (
	.clk(clk),
	.d(\Add2~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~2_combout ),
	.q(\processing_cnt[1]~q ),
	.prn(vcc));
defparam \processing_cnt[1] .is_wysiwyg = "true";
defparam \processing_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Add2~0 (
	.dataa(\processing_cnt[1]~q ),
	.datab(\processing_cnt[0]~q ),
	.datac(stg_valid_next),
	.datad(stg_sop_next),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout());
defparam \Add2~0 .lut_mask = 16'h6996;
defparam \Add2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add2~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\processing_cnt[2]~q ),
	.datad(\Add2~0_combout ),
	.cin(gnd),
	.combout(\Add2~1_combout ),
	.cout());
defparam \Add2~1 .lut_mask = 16'h0FF0;
defparam \Add2~1 .sum_lutc_input = "datac";

dffeas \processing_cnt[2] (
	.clk(clk),
	.d(\Add2~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\processing_cnt[2]~2_combout ),
	.q(\processing_cnt[2]~q ),
	.prn(vcc));
defparam \processing_cnt[2] .is_wysiwyg = "true";
defparam \processing_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \res~0 (
	.dataa(\processing_cnt[2]~q ),
	.datab(\processing_cnt[1]~q ),
	.datac(\processing_cnt[0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\res~0_combout ),
	.cout());
defparam \res~0 .lut_mask = 16'hFEFE;
defparam \res~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_bfi_1 (
	in_imag,
	in_real,
	out_stall_d,
	out_valid1,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	out_imag_2,
	out_real_2,
	out_inverse1,
	out_imag_3,
	out_real_3,
	out_imag_4,
	out_real_4,
	out_imag_5,
	out_real_5,
	out_imag_6,
	out_real_6,
	out_imag_7,
	out_real_7,
	out_imag_8,
	out_real_8,
	out_imag_9,
	out_real_9,
	out_eop1,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	out_sop_d_8,
	out_valid_d_8,
	out_inverse_d_8,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	[8:0] in_imag;
input 	[8:0] in_real;
input 	out_stall_d;
output 	out_valid1;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
output 	out_imag_2;
output 	out_real_2;
output 	out_inverse1;
output 	out_imag_3;
output 	out_real_3;
output 	out_imag_4;
output 	out_real_4;
output 	out_imag_5;
output 	out_real_5;
output 	out_imag_6;
output 	out_real_6;
output 	out_imag_7;
output 	out_real_7;
output 	out_imag_8;
output 	out_real_8;
output 	out_imag_9;
output 	out_real_9;
output 	out_eop1;
input 	fftpts_less_one_0;
input 	fftpts_less_one_1;
input 	fftpts_less_one_2;
input 	fftpts_less_one_3;
input 	out_sop_d_8;
input 	out_valid_d_8;
input 	out_inverse_d_8;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ;
wire \gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ;
wire \bf_control_inst|bf_counter_inst|control_s[0]~q ;
wire \bf_control_inst|out_valid~combout ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ;
wire \generate_delay_less_pipeline:in_imag_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ;
wire \generate_delay_less_pipeline:in_imag_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ;
wire \generate_delay_less_pipeline:in_imag_d[0]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ;
wire \generate_delay_less_pipeline:in_real_d[2]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ;
wire \generate_delay_less_pipeline:in_real_d[1]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ;
wire \generate_delay_less_pipeline:in_real_d[0]~q ;
wire \bf_control_inst|out_inverse~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ;
wire \generate_delay_less_pipeline:in_imag_d[3]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ;
wire \generate_delay_less_pipeline:in_real_d[3]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ;
wire \generate_delay_less_pipeline:in_imag_d[4]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ;
wire \generate_delay_less_pipeline:in_real_d[4]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ;
wire \generate_delay_less_pipeline:in_imag_d[5]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ;
wire \generate_delay_less_pipeline:in_real_d[5]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ;
wire \generate_delay_less_pipeline:in_imag_d[6]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ;
wire \generate_delay_less_pipeline:in_real_d[6]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ;
wire \generate_delay_less_pipeline:in_imag_d[7]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ;
wire \generate_delay_less_pipeline:in_real_d[7]~q ;
wire \generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ;
wire \generate_delay_less_pipeline:in_imag_d[8]~q ;
wire \generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ;
wire \generate_delay_less_pipeline:in_real_d[8]~q ;
wire \bf_control_inst|out_eop~q ;
wire \out_valid_d[0]~q ;
wire \out_valid_d[1]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ;
wire \s_sel_d[0]~q ;
wire \s_sel_d[1]~q ;
wire \out_imag~0_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ;
wire \out_real~0_combout ;
wire \out_inverse_d[0]~q ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ;
wire \out_imag~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ;
wire \out_real~1_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ;
wire \out_imag~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ;
wire \out_real~2_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ;
wire \out_imag~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ;
wire \out_real~3_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ;
wire \out_imag~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ;
wire \out_real~4_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ;
wire \out_imag~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ;
wire \out_real~5_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ;
wire \out_imag~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ;
wire \out_real~6_combout ;
wire \generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ;
wire \out_imag~7_combout ;
wire \generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ;
wire \out_real~7_combout ;
wire \out_eop_d[0]~q ;


ifft_8p_auk_dspip_r22sdf_bf_control_2 bf_control_inst(
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.enable(enable),
	.control_s_0(\bf_control_inst|bf_counter_inst|control_s[0]~q ),
	.out_valid1(\bf_control_inst|out_valid~combout ),
	.out_inverse1(\bf_control_inst|out_inverse~q ),
	.fftpts_less_one_0(fftpts_less_one_0),
	.fftpts_less_one_1(fftpts_less_one_1),
	.fftpts_less_one_2(fftpts_less_one_2),
	.fftpts_less_one_3(fftpts_less_one_3),
	.out_sop_d_8(out_sop_d_8),
	.out_valid_d_8(out_valid_d_8),
	.out_inverse_d_8(out_inverse_d_8),
	.out_eop1(\bf_control_inst|out_eop~q ),
	.clk(clk),
	.reset(reset));

ifft_8p_auk_dspip_r22sdf_addsub_10 \gen_fixedpt_adders:in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.generate_delay_less_pipelinein_imag_d2(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.generate_delay_less_pipelinein_imag_d1(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.generate_delay_less_pipelinein_imag_d0(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.generate_delay_less_pipelinein_imag_d3(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.generate_delay_less_pipelinein_imag_d4(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.generate_delay_less_pipelinein_imag_d5(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.generate_delay_less_pipelinein_imag_d6(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(\generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ),
	.generate_delay_less_pipelinein_imag_d7(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(\generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ),
	.generate_delay_less_pipelinein_imag_d8(\generate_delay_less_pipeline:in_imag_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_11 \gen_fixedpt_adders:in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d02(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.generate_delay_less_pipelinein_real_d2(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d01(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.generate_delay_less_pipelinein_real_d1(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d00(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.generate_delay_less_pipelinein_real_d0(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d03(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.generate_delay_less_pipelinein_real_d3(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d04(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.generate_delay_less_pipelinein_real_d4(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d05(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.generate_delay_less_pipelinein_real_d5(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d06(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.generate_delay_less_pipelinein_real_d6(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d07(\generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ),
	.generate_delay_less_pipelinein_real_d7(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d09(\generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ),
	.generate_delay_less_pipelinein_real_d8(\generate_delay_less_pipeline:in_real_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_8 \gen_fixedpt_adders:del_in_imag_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.generate_delay_less_pipelinein_imag_d2(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.generate_delay_less_pipelinein_imag_d1(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.generate_delay_less_pipelinein_imag_d0(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.generate_delay_less_pipelinein_imag_d3(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.generate_delay_less_pipelinein_imag_d4(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.generate_delay_less_pipelinein_imag_d5(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.generate_delay_less_pipelinein_imag_d6(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(\generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ),
	.generate_delay_less_pipelinein_imag_d7(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(\generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ),
	.generate_delay_less_pipelinein_imag_d8(\generate_delay_less_pipeline:in_imag_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_addsub_9 \gen_fixedpt_adders:del_in_real_comp_inst (
	.pipeline_dffe_2(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.pipeline_dffe_3(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.pipeline_dffe_4(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.pipeline_dffe_5(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.pipeline_dffe_6(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.pipeline_dffe_7(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.pipeline_dffe_8(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.pipeline_dffe_9(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.out_enable(enable),
	.generate_delay_less_pipelinedel_in_real_pl_d02(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.generate_delay_less_pipelinein_real_d2(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d01(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.generate_delay_less_pipelinein_real_d1(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d00(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.generate_delay_less_pipelinein_real_d0(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d03(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.generate_delay_less_pipelinein_real_d3(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d04(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.generate_delay_less_pipelinein_real_d4(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d05(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.generate_delay_less_pipelinein_real_d5(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d06(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.generate_delay_less_pipelinein_real_d6(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d07(\generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ),
	.generate_delay_less_pipelinein_real_d7(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.generate_delay_less_pipelinedel_in_real_pl_d09(\generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ),
	.generate_delay_less_pipelinein_real_d8(\generate_delay_less_pipeline:in_real_d[8]~q ),
	.clk(clk),
	.reset_n(reset));

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[2] (
	.clk(clk),
	.d(in_imag[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[1] (
	.clk(clk),
	.d(in_imag[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[0] (
	.clk(clk),
	.d(in_imag[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][2] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][2] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[2] (
	.clk(clk),
	.d(in_real[2]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[2] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][1] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][1] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[1] (
	.clk(clk),
	.d(in_real[1]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[1]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[1] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][0] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][0] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[0] (
	.clk(clk),
	.d(in_real[0]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[0]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[0] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[3] (
	.clk(clk),
	.d(in_imag[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][3] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][3] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[3] (
	.clk(clk),
	.d(in_real[3]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[3] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[4] (
	.clk(clk),
	.d(in_imag[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][4] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][4] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[4] (
	.clk(clk),
	.d(in_real[4]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[4] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[5] (
	.clk(clk),
	.d(in_imag[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][5] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][5] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[5] (
	.clk(clk),
	.d(in_real[5]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[5] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[6] (
	.clk(clk),
	.d(in_imag[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][6] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][6] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[6] (
	.clk(clk),
	.d(in_real[6]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[6] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[7] (
	.clk(clk),
	.d(in_imag[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][7] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][7] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[7] (
	.clk(clk),
	.d(in_real[7]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[7] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_imag_d[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_imag_pl_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_imag_pl_d[0][9] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_imag_d[8] (
	.clk(clk),
	.d(in_imag[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_imag_d[8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_imag_d[8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_imag_d[8] .power_up = "low";

dffeas \generate_delay_less_pipeline:del_in_real_pl_d[0][9] (
	.clk(clk),
	.d(\generate_delay_less_pipeline:in_real_d[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:del_in_real_pl_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:del_in_real_pl_d[0][9] .power_up = "low";

dffeas \generate_delay_less_pipeline:in_real_d[8] (
	.clk(clk),
	.d(in_real[8]),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:in_real_d[8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:in_real_d[8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:in_real_d[8] .power_up = "low";

dffeas out_valid(
	.clk(clk),
	.d(\out_valid_d[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_valid1),
	.prn(vcc));
defparam out_valid.is_wysiwyg = "true";
defparam out_valid.power_up = "low";

dffeas \out_imag[2] (
	.clk(clk),
	.d(\out_imag~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_2),
	.prn(vcc));
defparam \out_imag[2] .is_wysiwyg = "true";
defparam \out_imag[2] .power_up = "low";

dffeas \out_real[2] (
	.clk(clk),
	.d(\out_real~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_2),
	.prn(vcc));
defparam \out_real[2] .is_wysiwyg = "true";
defparam \out_real[2] .power_up = "low";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

dffeas \out_imag[3] (
	.clk(clk),
	.d(\out_imag~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_3),
	.prn(vcc));
defparam \out_imag[3] .is_wysiwyg = "true";
defparam \out_imag[3] .power_up = "low";

dffeas \out_real[3] (
	.clk(clk),
	.d(\out_real~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_3),
	.prn(vcc));
defparam \out_real[3] .is_wysiwyg = "true";
defparam \out_real[3] .power_up = "low";

dffeas \out_imag[4] (
	.clk(clk),
	.d(\out_imag~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_4),
	.prn(vcc));
defparam \out_imag[4] .is_wysiwyg = "true";
defparam \out_imag[4] .power_up = "low";

dffeas \out_real[4] (
	.clk(clk),
	.d(\out_real~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_4),
	.prn(vcc));
defparam \out_real[4] .is_wysiwyg = "true";
defparam \out_real[4] .power_up = "low";

dffeas \out_imag[5] (
	.clk(clk),
	.d(\out_imag~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_5),
	.prn(vcc));
defparam \out_imag[5] .is_wysiwyg = "true";
defparam \out_imag[5] .power_up = "low";

dffeas \out_real[5] (
	.clk(clk),
	.d(\out_real~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_5),
	.prn(vcc));
defparam \out_real[5] .is_wysiwyg = "true";
defparam \out_real[5] .power_up = "low";

dffeas \out_imag[6] (
	.clk(clk),
	.d(\out_imag~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_6),
	.prn(vcc));
defparam \out_imag[6] .is_wysiwyg = "true";
defparam \out_imag[6] .power_up = "low";

dffeas \out_real[6] (
	.clk(clk),
	.d(\out_real~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_6),
	.prn(vcc));
defparam \out_real[6] .is_wysiwyg = "true";
defparam \out_real[6] .power_up = "low";

dffeas \out_imag[7] (
	.clk(clk),
	.d(\out_imag~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_7),
	.prn(vcc));
defparam \out_imag[7] .is_wysiwyg = "true";
defparam \out_imag[7] .power_up = "low";

dffeas \out_real[7] (
	.clk(clk),
	.d(\out_real~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_7),
	.prn(vcc));
defparam \out_real[7] .is_wysiwyg = "true";
defparam \out_real[7] .power_up = "low";

dffeas \out_imag[8] (
	.clk(clk),
	.d(\out_imag~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_8),
	.prn(vcc));
defparam \out_imag[8] .is_wysiwyg = "true";
defparam \out_imag[8] .power_up = "low";

dffeas \out_real[8] (
	.clk(clk),
	.d(\out_real~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_8),
	.prn(vcc));
defparam \out_real[8] .is_wysiwyg = "true";
defparam \out_real[8] .power_up = "low";

dffeas \out_imag[9] (
	.clk(clk),
	.d(\out_imag~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_imag_9),
	.prn(vcc));
defparam \out_imag[9] .is_wysiwyg = "true";
defparam \out_imag[9] .power_up = "low";

dffeas \out_real[9] (
	.clk(clk),
	.d(\out_real~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_real_9),
	.prn(vcc));
defparam \out_real[9] .is_wysiwyg = "true";
defparam \out_real[9] .power_up = "low";

dffeas out_eop(
	.clk(clk),
	.d(\out_eop_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_eop1),
	.prn(vcc));
defparam out_eop.is_wysiwyg = "true";
defparam out_eop.power_up = "low";

dffeas \out_valid_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_valid~combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[0]~q ),
	.prn(vcc));
defparam \out_valid_d[0] .is_wysiwyg = "true";
defparam \out_valid_d[0] .power_up = "low";

dffeas \out_valid_d[1] (
	.clk(clk),
	.d(\out_valid_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_valid_d[1]~q ),
	.prn(vcc));
defparam \out_valid_d[1] .is_wysiwyg = "true";
defparam \out_valid_d[1] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][2] .power_up = "low";

dffeas \s_sel_d[0] (
	.clk(clk),
	.d(\bf_control_inst|bf_counter_inst|control_s[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[0]~q ),
	.prn(vcc));
defparam \s_sel_d[0] .is_wysiwyg = "true";
defparam \s_sel_d[0] .power_up = "low";

dffeas \s_sel_d[1] (
	.clk(clk),
	.d(\s_sel_d[0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\s_sel_d[1]~q ),
	.prn(vcc));
defparam \s_sel_d[1] .is_wysiwyg = "true";
defparam \s_sel_d[1] .power_up = "low";

cycloneiv_lcell_comb \out_imag~0 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][2]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~0_combout ),
	.cout());
defparam \out_imag~0 .lut_mask = 16'hAACC;
defparam \out_imag~0 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][2] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][2] .power_up = "low";

cycloneiv_lcell_comb \out_real~0 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][2]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~0_combout ),
	.cout());
defparam \out_real~0 .lut_mask = 16'hAACC;
defparam \out_real~0 .sum_lutc_input = "datac";

dffeas \out_inverse_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_inverse~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_inverse_d[0]~q ),
	.prn(vcc));
defparam \out_inverse_d[0] .is_wysiwyg = "true";
defparam \out_inverse_d[0] .power_up = "low";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \out_imag~1 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][3]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~1_combout ),
	.cout());
defparam \out_imag~1 .lut_mask = 16'hAACC;
defparam \out_imag~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][3] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][3] .power_up = "low";

cycloneiv_lcell_comb \out_real~1 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][3]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~1_combout ),
	.cout());
defparam \out_real~1 .lut_mask = 16'hAACC;
defparam \out_real~1 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \out_imag~2 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][4]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~2_combout ),
	.cout());
defparam \out_imag~2 .lut_mask = 16'hAACC;
defparam \out_imag~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][4] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][4] .power_up = "low";

cycloneiv_lcell_comb \out_real~2 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][4]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~2_combout ),
	.cout());
defparam \out_real~2 .lut_mask = 16'hAACC;
defparam \out_real~2 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \out_imag~3 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][5]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~3_combout ),
	.cout());
defparam \out_imag~3 .lut_mask = 16'hAACC;
defparam \out_imag~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][5] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][5] .power_up = "low";

cycloneiv_lcell_comb \out_real~3 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][5]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~3_combout ),
	.cout());
defparam \out_real~3 .lut_mask = 16'hAACC;
defparam \out_real~3 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \out_imag~4 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][6]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~4_combout ),
	.cout());
defparam \out_imag~4 .lut_mask = 16'hAACC;
defparam \out_imag~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][6] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][6] .power_up = "low";

cycloneiv_lcell_comb \out_real~4 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][6]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~4_combout ),
	.cout());
defparam \out_real~4 .lut_mask = 16'hAACC;
defparam \out_real~4 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][7] .power_up = "low";

cycloneiv_lcell_comb \out_imag~5 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][7]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~5_combout ),
	.cout());
defparam \out_imag~5 .lut_mask = 16'hAACC;
defparam \out_imag~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][7] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][7] .power_up = "low";

cycloneiv_lcell_comb \out_real~5 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][7]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~5_combout ),
	.cout());
defparam \out_real~5 .lut_mask = 16'hAACC;
defparam \out_real~5 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][8] .power_up = "low";

cycloneiv_lcell_comb \out_imag~6 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][8]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~6_combout ),
	.cout());
defparam \out_imag~6 .lut_mask = 16'hAACC;
defparam \out_imag~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][8] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][8] .power_up = "low";

cycloneiv_lcell_comb \out_real~6 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][8]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~6_combout ),
	.cout());
defparam \out_real~6 .lut_mask = 16'hAACC;
defparam \out_real~6 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_imag_d[0][9] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_imag_d[0][9] .power_up = "low";

cycloneiv_lcell_comb \out_imag~7 (
	.dataa(\gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_imag_d[0][9]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_imag~7_combout ),
	.cout());
defparam \out_imag~7 .lut_mask = 16'hAACC;
defparam \out_imag~7 .sum_lutc_input = "datac";

dffeas \generate_delay_less_pipeline:adder2_out_real_d[0][9] (
	.clk(clk),
	.d(\gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ),
	.prn(vcc));
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][9] .is_wysiwyg = "true";
defparam \generate_delay_less_pipeline:adder2_out_real_d[0][9] .power_up = "low";

cycloneiv_lcell_comb \out_real~7 (
	.dataa(\gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~q ),
	.datab(\generate_delay_less_pipeline:adder2_out_real_d[0][9]~q ),
	.datac(gnd),
	.datad(\s_sel_d[1]~q ),
	.cin(gnd),
	.combout(\out_real~7_combout ),
	.cout());
defparam \out_real~7 .lut_mask = 16'hAACC;
defparam \out_real~7 .sum_lutc_input = "datac";

dffeas \out_eop_d[0] (
	.clk(clk),
	.d(\bf_control_inst|out_eop~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\out_eop_d[0]~q ),
	.prn(vcc));
defparam \out_eop_d[0] .is_wysiwyg = "true";
defparam \out_eop_d[0] .power_up = "low";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_8 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_9 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.generate_delay_less_pipelinein_imag_d8(generate_delay_less_pipelinein_imag_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_4 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.generate_delay_less_pipelinein_imag_d8(generate_delay_less_pipelinein_imag_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_4 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.datab(generate_delay_less_pipelinein_imag_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00EE;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.datab(generate_delay_less_pipelinein_imag_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h007F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.datab(generate_delay_less_pipelinein_imag_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.datab(generate_delay_less_pipelinein_imag_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.datab(generate_delay_less_pipelinein_imag_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.datab(generate_delay_less_pipelinein_imag_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.datab(generate_delay_less_pipelinein_imag_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.datab(generate_delay_less_pipelinein_imag_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.datab(generate_delay_less_pipelinein_imag_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_9 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_10 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d02(generate_delay_less_pipelinedel_in_real_pl_d02),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d01(generate_delay_less_pipelinedel_in_real_pl_d01),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d00(generate_delay_less_pipelinedel_in_real_pl_d00),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d03(generate_delay_less_pipelinedel_in_real_pl_d03),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d04(generate_delay_less_pipelinedel_in_real_pl_d04),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d05(generate_delay_less_pipelinedel_in_real_pl_d05),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d06(generate_delay_less_pipelinedel_in_real_pl_d06),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d07(generate_delay_less_pipelinedel_in_real_pl_d07),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d09(generate_delay_less_pipelinedel_in_real_pl_d09),
	.generate_delay_less_pipelinein_real_d8(generate_delay_less_pipelinein_real_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_5 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d02(generate_delay_less_pipelinedel_in_real_pl_d02),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d01(generate_delay_less_pipelinedel_in_real_pl_d01),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d00(generate_delay_less_pipelinedel_in_real_pl_d00),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d03(generate_delay_less_pipelinedel_in_real_pl_d03),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d04(generate_delay_less_pipelinedel_in_real_pl_d04),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d05(generate_delay_less_pipelinedel_in_real_pl_d05),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d06(generate_delay_less_pipelinedel_in_real_pl_d06),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d07(generate_delay_less_pipelinedel_in_real_pl_d07),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d09(generate_delay_less_pipelinedel_in_real_pl_d09),
	.generate_delay_less_pipelinein_real_d8(generate_delay_less_pipelinein_real_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_5 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d00),
	.datab(generate_delay_less_pipelinein_real_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00EE;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d01),
	.datab(generate_delay_less_pipelinein_real_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h007F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d02),
	.datab(generate_delay_less_pipelinein_real_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d03),
	.datab(generate_delay_less_pipelinein_real_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d04),
	.datab(generate_delay_less_pipelinein_real_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d05),
	.datab(generate_delay_less_pipelinein_real_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d06),
	.datab(generate_delay_less_pipelinein_real_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d07),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h967F;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d09),
	.datab(generate_delay_less_pipelinein_real_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96EF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d09),
	.datab(generate_delay_less_pipelinein_real_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:del_in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_10 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_11 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.generate_delay_less_pipelinein_imag_d8(generate_delay_less_pipelinein_imag_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_6 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_imag_pl_d02(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.generate_delay_less_pipelinein_imag_d2(generate_delay_less_pipelinein_imag_d2),
	.generate_delay_less_pipelinedel_in_imag_pl_d01(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.generate_delay_less_pipelinein_imag_d1(generate_delay_less_pipelinein_imag_d1),
	.generate_delay_less_pipelinedel_in_imag_pl_d00(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.generate_delay_less_pipelinein_imag_d0(generate_delay_less_pipelinein_imag_d0),
	.generate_delay_less_pipelinedel_in_imag_pl_d03(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.generate_delay_less_pipelinein_imag_d3(generate_delay_less_pipelinein_imag_d3),
	.generate_delay_less_pipelinedel_in_imag_pl_d04(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.generate_delay_less_pipelinein_imag_d4(generate_delay_less_pipelinein_imag_d4),
	.generate_delay_less_pipelinedel_in_imag_pl_d05(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.generate_delay_less_pipelinein_imag_d5(generate_delay_less_pipelinein_imag_d5),
	.generate_delay_less_pipelinedel_in_imag_pl_d06(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.generate_delay_less_pipelinein_imag_d6(generate_delay_less_pipelinein_imag_d6),
	.generate_delay_less_pipelinedel_in_imag_pl_d07(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.generate_delay_less_pipelinein_imag_d7(generate_delay_less_pipelinein_imag_d7),
	.generate_delay_less_pipelinedel_in_imag_pl_d09(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.generate_delay_less_pipelinein_imag_d8(generate_delay_less_pipelinein_imag_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_6 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_imag_pl_d02,
	generate_delay_less_pipelinein_imag_d2,
	generate_delay_less_pipelinedel_in_imag_pl_d01,
	generate_delay_less_pipelinein_imag_d1,
	generate_delay_less_pipelinedel_in_imag_pl_d00,
	generate_delay_less_pipelinein_imag_d0,
	generate_delay_less_pipelinedel_in_imag_pl_d03,
	generate_delay_less_pipelinein_imag_d3,
	generate_delay_less_pipelinedel_in_imag_pl_d04,
	generate_delay_less_pipelinein_imag_d4,
	generate_delay_less_pipelinedel_in_imag_pl_d05,
	generate_delay_less_pipelinein_imag_d5,
	generate_delay_less_pipelinedel_in_imag_pl_d06,
	generate_delay_less_pipelinein_imag_d6,
	generate_delay_less_pipelinedel_in_imag_pl_d07,
	generate_delay_less_pipelinein_imag_d7,
	generate_delay_less_pipelinedel_in_imag_pl_d09,
	generate_delay_less_pipelinein_imag_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_imag_pl_d02;
input 	generate_delay_less_pipelinein_imag_d2;
input 	generate_delay_less_pipelinedel_in_imag_pl_d01;
input 	generate_delay_less_pipelinein_imag_d1;
input 	generate_delay_less_pipelinedel_in_imag_pl_d00;
input 	generate_delay_less_pipelinein_imag_d0;
input 	generate_delay_less_pipelinedel_in_imag_pl_d03;
input 	generate_delay_less_pipelinein_imag_d3;
input 	generate_delay_less_pipelinedel_in_imag_pl_d04;
input 	generate_delay_less_pipelinein_imag_d4;
input 	generate_delay_less_pipelinedel_in_imag_pl_d05;
input 	generate_delay_less_pipelinein_imag_d5;
input 	generate_delay_less_pipelinedel_in_imag_pl_d06;
input 	generate_delay_less_pipelinein_imag_d6;
input 	generate_delay_less_pipelinedel_in_imag_pl_d07;
input 	generate_delay_less_pipelinein_imag_d7;
input 	generate_delay_less_pipelinedel_in_imag_pl_d09;
input 	generate_delay_less_pipelinein_imag_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d00),
	.datab(generate_delay_less_pipelinein_imag_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00BB;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d01),
	.datab(generate_delay_less_pipelinein_imag_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h00DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d02),
	.datab(generate_delay_less_pipelinein_imag_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d03),
	.datab(generate_delay_less_pipelinein_imag_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d04),
	.datab(generate_delay_less_pipelinein_imag_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d05),
	.datab(generate_delay_less_pipelinein_imag_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d06),
	.datab(generate_delay_less_pipelinein_imag_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d07),
	.datab(generate_delay_less_pipelinein_imag_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.datab(generate_delay_less_pipelinein_imag_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_imag_pl_d09),
	.datab(generate_delay_less_pipelinein_imag_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_imag_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_addsub_11 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	out_enable,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	out_enable;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_LPM_ADD_SUB_12 \gen_pipeline:lpm_add_sub_component (
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(out_enable),
	.generate_delay_less_pipelinedel_in_real_pl_d02(generate_delay_less_pipelinedel_in_real_pl_d02),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d01(generate_delay_less_pipelinedel_in_real_pl_d01),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d00(generate_delay_less_pipelinedel_in_real_pl_d00),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d03(generate_delay_less_pipelinedel_in_real_pl_d03),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d04(generate_delay_less_pipelinedel_in_real_pl_d04),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d05(generate_delay_less_pipelinedel_in_real_pl_d05),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d06(generate_delay_less_pipelinedel_in_real_pl_d06),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d07(generate_delay_less_pipelinedel_in_real_pl_d07),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d09(generate_delay_less_pipelinedel_in_real_pl_d09),
	.generate_delay_less_pipelinein_real_d8(generate_delay_less_pipelinein_real_d8),
	.clock(clk),
	.reset_n(reset_n));

endmodule

module ifft_8p_LPM_ADD_SUB_12 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_add_sub_4ij_7 auto_generated(
	.pipeline_dffe_2(pipeline_dffe_2),
	.pipeline_dffe_3(pipeline_dffe_3),
	.pipeline_dffe_4(pipeline_dffe_4),
	.pipeline_dffe_5(pipeline_dffe_5),
	.pipeline_dffe_6(pipeline_dffe_6),
	.pipeline_dffe_7(pipeline_dffe_7),
	.pipeline_dffe_8(pipeline_dffe_8),
	.pipeline_dffe_9(pipeline_dffe_9),
	.clken(clken),
	.generate_delay_less_pipelinedel_in_real_pl_d02(generate_delay_less_pipelinedel_in_real_pl_d02),
	.generate_delay_less_pipelinein_real_d2(generate_delay_less_pipelinein_real_d2),
	.generate_delay_less_pipelinedel_in_real_pl_d01(generate_delay_less_pipelinedel_in_real_pl_d01),
	.generate_delay_less_pipelinein_real_d1(generate_delay_less_pipelinein_real_d1),
	.generate_delay_less_pipelinedel_in_real_pl_d00(generate_delay_less_pipelinedel_in_real_pl_d00),
	.generate_delay_less_pipelinein_real_d0(generate_delay_less_pipelinein_real_d0),
	.generate_delay_less_pipelinedel_in_real_pl_d03(generate_delay_less_pipelinedel_in_real_pl_d03),
	.generate_delay_less_pipelinein_real_d3(generate_delay_less_pipelinein_real_d3),
	.generate_delay_less_pipelinedel_in_real_pl_d04(generate_delay_less_pipelinedel_in_real_pl_d04),
	.generate_delay_less_pipelinein_real_d4(generate_delay_less_pipelinein_real_d4),
	.generate_delay_less_pipelinedel_in_real_pl_d05(generate_delay_less_pipelinedel_in_real_pl_d05),
	.generate_delay_less_pipelinein_real_d5(generate_delay_less_pipelinein_real_d5),
	.generate_delay_less_pipelinedel_in_real_pl_d06(generate_delay_less_pipelinedel_in_real_pl_d06),
	.generate_delay_less_pipelinein_real_d6(generate_delay_less_pipelinein_real_d6),
	.generate_delay_less_pipelinedel_in_real_pl_d07(generate_delay_less_pipelinedel_in_real_pl_d07),
	.generate_delay_less_pipelinein_real_d7(generate_delay_less_pipelinein_real_d7),
	.generate_delay_less_pipelinedel_in_real_pl_d09(generate_delay_less_pipelinedel_in_real_pl_d09),
	.generate_delay_less_pipelinein_real_d8(generate_delay_less_pipelinein_real_d8),
	.clock(clock),
	.reset_n(reset_n));

endmodule

module ifft_8p_add_sub_4ij_7 (
	pipeline_dffe_2,
	pipeline_dffe_3,
	pipeline_dffe_4,
	pipeline_dffe_5,
	pipeline_dffe_6,
	pipeline_dffe_7,
	pipeline_dffe_8,
	pipeline_dffe_9,
	clken,
	generate_delay_less_pipelinedel_in_real_pl_d02,
	generate_delay_less_pipelinein_real_d2,
	generate_delay_less_pipelinedel_in_real_pl_d01,
	generate_delay_less_pipelinein_real_d1,
	generate_delay_less_pipelinedel_in_real_pl_d00,
	generate_delay_less_pipelinein_real_d0,
	generate_delay_less_pipelinedel_in_real_pl_d03,
	generate_delay_less_pipelinein_real_d3,
	generate_delay_less_pipelinedel_in_real_pl_d04,
	generate_delay_less_pipelinein_real_d4,
	generate_delay_less_pipelinedel_in_real_pl_d05,
	generate_delay_less_pipelinein_real_d5,
	generate_delay_less_pipelinedel_in_real_pl_d06,
	generate_delay_less_pipelinein_real_d6,
	generate_delay_less_pipelinedel_in_real_pl_d07,
	generate_delay_less_pipelinein_real_d7,
	generate_delay_less_pipelinedel_in_real_pl_d09,
	generate_delay_less_pipelinein_real_d8,
	clock,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	pipeline_dffe_2;
output 	pipeline_dffe_3;
output 	pipeline_dffe_4;
output 	pipeline_dffe_5;
output 	pipeline_dffe_6;
output 	pipeline_dffe_7;
output 	pipeline_dffe_8;
output 	pipeline_dffe_9;
input 	clken;
input 	generate_delay_less_pipelinedel_in_real_pl_d02;
input 	generate_delay_less_pipelinein_real_d2;
input 	generate_delay_less_pipelinedel_in_real_pl_d01;
input 	generate_delay_less_pipelinein_real_d1;
input 	generate_delay_less_pipelinedel_in_real_pl_d00;
input 	generate_delay_less_pipelinein_real_d0;
input 	generate_delay_less_pipelinedel_in_real_pl_d03;
input 	generate_delay_less_pipelinein_real_d3;
input 	generate_delay_less_pipelinedel_in_real_pl_d04;
input 	generate_delay_less_pipelinein_real_d4;
input 	generate_delay_less_pipelinedel_in_real_pl_d05;
input 	generate_delay_less_pipelinein_real_d5;
input 	generate_delay_less_pipelinedel_in_real_pl_d06;
input 	generate_delay_less_pipelinein_real_d6;
input 	generate_delay_less_pipelinedel_in_real_pl_d07;
input 	generate_delay_less_pipelinein_real_d7;
input 	generate_delay_less_pipelinedel_in_real_pl_d09;
input 	generate_delay_less_pipelinein_real_d8;
input 	clock;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ;
wire \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ;


dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_2),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_3),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_4),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_5),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_6),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_7),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_8),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8] .power_up = "low";

dffeas \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] (
	.clk(clock),
	.d(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(clken),
	.q(pipeline_dffe_9),
	.prn(vcc));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .is_wysiwyg = "true";
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9] .power_up = "low";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d00),
	.datab(generate_delay_less_pipelinein_real_d0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .lut_mask = 16'h00BB;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d01),
	.datab(generate_delay_less_pipelinein_real_d1),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~9_cout ),
	.combout(),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .lut_mask = 16'h00DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d02),
	.datab(generate_delay_less_pipelinein_real_d2),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~11_cout ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d03),
	.datab(generate_delay_less_pipelinein_real_d3),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[2]~13 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d04),
	.datab(generate_delay_less_pipelinein_real_d4),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[3]~15 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d05),
	.datab(generate_delay_less_pipelinein_real_d5),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[4]~17 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d06),
	.datab(generate_delay_less_pipelinein_real_d6),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[5]~19 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d07),
	.datab(generate_delay_less_pipelinein_real_d7),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[6]~21 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .lut_mask = 16'h96DF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d09),
	.datab(generate_delay_less_pipelinein_real_d8),
	.datac(gnd),
	.datad(vcc),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[7]~23 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24_combout ),
	.cout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ));
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .lut_mask = 16'h96BF;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 (
	.dataa(generate_delay_less_pipelinedel_in_real_pl_d09),
	.datab(generate_delay_less_pipelinein_real_d8),
	.datac(gnd),
	.datad(gnd),
	.cin(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[8]~25 ),
	.combout(\fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26_combout ),
	.cout());
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .lut_mask = 16'h9696;
defparam \fft_ii_0|auk_dspip_r22sdf_top_inst|r22sdf_core_inst|gen_natural_order_core:gen_stages:1:r22_stage|gen_bfi:gen_bfi_only:bfi_inst|gen_fixedpt_adders:in_real_comp_inst|gen_pipeline:lpm_add_sub_component|auto_generated|pipeline_dffe[9]~26 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_bf_control_2 (
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	enable,
	control_s_0,
	out_valid1,
	out_inverse1,
	fftpts_less_one_0,
	fftpts_less_one_1,
	fftpts_less_one_2,
	fftpts_less_one_3,
	out_sop_d_8,
	out_valid_d_8,
	out_inverse_d_8,
	out_eop1,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	enable;
output 	control_s_0;
output 	out_valid1;
output 	out_inverse1;
input 	fftpts_less_one_0;
input 	fftpts_less_one_1;
input 	fftpts_less_one_2;
input 	fftpts_less_one_3;
input 	out_sop_d_8;
input 	out_valid_d_8;
input 	out_inverse_d_8;
output 	out_eop1;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \bf_counter_inst|counter_p~0_combout ;
wire \Add3~1_combout ;
wire \in_cnt~2_combout ;
wire \in_cnt[2]~q ;
wire \Add3~0_combout ;
wire \in_cnt~1_combout ;
wire \in_cnt[3]~q ;
wire \Equal0~1_combout ;
wire \in_cnt~3_combout ;
wire \in_cnt[1]~q ;
wire \Equal0~0_combout ;
wire \in_cnt~0_combout ;
wire \in_cnt[0]~q ;
wire \gen_out_cnt_p~0_combout ;
wire \gen_out_cnt_p~1_combout ;
wire \Add4~1_combout ;
wire \out_cnt[2]~7_combout ;
wire \out_cnt[2]~q ;
wire \Add4~0_combout ;
wire \out_cnt[3]~6_combout ;
wire \out_cnt[3]~q ;
wire \Equal2~1_combout ;
wire \out_cnt[3]~3_combout ;
wire \out_cnt[0]~5_combout ;
wire \out_cnt[0]~q ;
wire \out_cnt[3]~0_combout ;
wire \out_cnt[3]~1_combout ;
wire \out_cnt[3]~2_combout ;
wire \out_cnt[1]~4_combout ;
wire \out_cnt[1]~q ;
wire \Equal2~0_combout ;
wire \shift~0_combout ;
wire \shift~q ;
wire \out_inverse~0_combout ;


ifft_8p_auk_dspip_r22sdf_counter_2 bf_counter_inst(
	.out_stall_d(out_stall_d),
	.curr_pwr_2_s(curr_pwr_2_s),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.control_s_0(control_s_0),
	.out_sop_d_8(out_sop_d_8),
	.out_valid_d_8(out_valid_d_8),
	.counter_p(\bf_counter_inst|counter_p~0_combout ),
	.clk(clk),
	.reset(reset));

cycloneiv_lcell_comb out_valid(
	.dataa(\shift~q ),
	.datab(control_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(out_valid1),
	.cout());
defparam out_valid.lut_mask = 16'hEEEE;
defparam out_valid.sum_lutc_input = "datac";

dffeas out_inverse(
	.clk(clk),
	.d(\out_inverse~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(out_inverse1),
	.prn(vcc));
defparam out_inverse.is_wysiwyg = "true";
defparam out_inverse.power_up = "low";

dffeas out_eop(
	.clk(clk),
	.d(\out_cnt[3]~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(out_eop1),
	.prn(vcc));
defparam out_eop.is_wysiwyg = "true";
defparam out_eop.power_up = "low";

cycloneiv_lcell_comb \Add3~1 (
	.dataa(gnd),
	.datab(\in_cnt[2]~q ),
	.datac(\in_cnt[0]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add3~1_combout ),
	.cout());
defparam \Add3~1 .lut_mask = 16'hC33C;
defparam \Add3~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~2 (
	.dataa(\Add3~1_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~2_combout ),
	.cout());
defparam \in_cnt~2 .lut_mask = 16'hAFFF;
defparam \in_cnt~2 .sum_lutc_input = "datac";

dffeas \in_cnt[2] (
	.clk(clk),
	.d(\in_cnt~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[2]~q ),
	.prn(vcc));
defparam \in_cnt[2] .is_wysiwyg = "true";
defparam \in_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Add3~0 (
	.dataa(\in_cnt[3]~q ),
	.datab(\in_cnt[0]~q ),
	.datac(\in_cnt[2]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout());
defparam \Add3~0 .lut_mask = 16'h6996;
defparam \Add3~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~1 (
	.dataa(\Add3~0_combout ),
	.datab(gnd),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~1_combout ),
	.cout());
defparam \in_cnt~1 .lut_mask = 16'hAFFF;
defparam \in_cnt~1 .sum_lutc_input = "datac";

dffeas \in_cnt[3] (
	.clk(clk),
	.d(\in_cnt~1_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[3]~q ),
	.prn(vcc));
defparam \in_cnt[3] .is_wysiwyg = "true";
defparam \in_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \Equal0~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\in_cnt[3]~q ),
	.datad(\in_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal0~1_combout ),
	.cout());
defparam \Equal0~1 .lut_mask = 16'h6996;
defparam \Equal0~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~3 (
	.dataa(\in_cnt[0]~q ),
	.datab(\in_cnt[1]~q ),
	.datac(\Equal0~0_combout ),
	.datad(\Equal0~1_combout ),
	.cin(gnd),
	.combout(\in_cnt~3_combout ),
	.cout());
defparam \in_cnt~3 .lut_mask = 16'h6FFF;
defparam \in_cnt~3 .sum_lutc_input = "datac";

dffeas \in_cnt[1] (
	.clk(clk),
	.d(\in_cnt~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[1]~q ),
	.prn(vcc));
defparam \in_cnt[1] .is_wysiwyg = "true";
defparam \in_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal0~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\in_cnt[1]~q ),
	.datad(\in_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
defparam \Equal0~0 .lut_mask = 16'h6996;
defparam \Equal0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_cnt~0 (
	.dataa(\in_cnt[0]~q ),
	.datab(\Equal0~0_combout ),
	.datac(\Equal0~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_cnt~0_combout ),
	.cout());
defparam \in_cnt~0 .lut_mask = 16'h7F7F;
defparam \in_cnt~0 .sum_lutc_input = "datac";

dffeas \in_cnt[0] (
	.clk(clk),
	.d(\in_cnt~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\bf_counter_inst|counter_p~0_combout ),
	.q(\in_cnt[0]~q ),
	.prn(vcc));
defparam \in_cnt[0] .is_wysiwyg = "true";
defparam \in_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \gen_out_cnt_p~0 (
	.dataa(curr_pwr_2_s),
	.datab(\in_cnt[3]~q ),
	.datac(\in_cnt[2]~q ),
	.datad(\in_cnt[1]~q ),
	.cin(gnd),
	.combout(\gen_out_cnt_p~0_combout ),
	.cout());
defparam \gen_out_cnt_p~0 .lut_mask = 16'hBFFF;
defparam \gen_out_cnt_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \gen_out_cnt_p~1 (
	.dataa(\in_cnt[0]~q ),
	.datab(\gen_out_cnt_p~0_combout ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\gen_out_cnt_p~1_combout ),
	.cout());
defparam \gen_out_cnt_p~1 .lut_mask = 16'hEEEE;
defparam \gen_out_cnt_p~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~1 (
	.dataa(gnd),
	.datab(\out_cnt[2]~q ),
	.datac(\out_cnt[0]~q ),
	.datad(\out_cnt[1]~q ),
	.cin(gnd),
	.combout(\Add4~1_combout ),
	.cout());
defparam \Add4~1 .lut_mask = 16'hC33C;
defparam \Add4~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[2]~7 (
	.dataa(\out_cnt[2]~q ),
	.datab(\out_cnt[3]~3_combout ),
	.datac(\Add4~1_combout ),
	.datad(\out_cnt[3]~2_combout ),
	.cin(gnd),
	.combout(\out_cnt[2]~7_combout ),
	.cout());
defparam \out_cnt[2]~7 .lut_mask = 16'hBBF3;
defparam \out_cnt[2]~7 .sum_lutc_input = "datac";

dffeas \out_cnt[2] (
	.clk(clk),
	.d(\out_cnt[2]~7_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[2]~q ),
	.prn(vcc));
defparam \out_cnt[2] .is_wysiwyg = "true";
defparam \out_cnt[2] .power_up = "low";

cycloneiv_lcell_comb \Add4~0 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[0]~q ),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout());
defparam \Add4~0 .lut_mask = 16'h6996;
defparam \Add4~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~6 (
	.dataa(\out_cnt[3]~q ),
	.datab(\out_cnt[3]~3_combout ),
	.datac(\Add4~0_combout ),
	.datad(\out_cnt[3]~2_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~6_combout ),
	.cout());
defparam \out_cnt[3]~6 .lut_mask = 16'hBBF3;
defparam \out_cnt[3]~6 .sum_lutc_input = "datac";

dffeas \out_cnt[3] (
	.clk(clk),
	.d(\out_cnt[3]~6_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[3]~q ),
	.prn(vcc));
defparam \out_cnt[3] .is_wysiwyg = "true";
defparam \out_cnt[3] .power_up = "low";

cycloneiv_lcell_comb \Equal2~1 (
	.dataa(fftpts_less_one_2),
	.datab(fftpts_less_one_3),
	.datac(\out_cnt[3]~q ),
	.datad(\out_cnt[2]~q ),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
defparam \Equal2~1 .lut_mask = 16'h6996;
defparam \Equal2~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~3 (
	.dataa(\in_cnt[0]~q ),
	.datab(\gen_out_cnt_p~0_combout ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~3_combout ),
	.cout());
defparam \out_cnt[3]~3 .lut_mask = 16'hFFF7;
defparam \out_cnt[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[0]~5 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(\out_cnt[3]~3_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_cnt[0]~5_combout ),
	.cout());
defparam \out_cnt[0]~5 .lut_mask = 16'h6F6F;
defparam \out_cnt[0]~5 .sum_lutc_input = "datac";

dffeas \out_cnt[0] (
	.clk(clk),
	.d(\out_cnt[0]~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[0]~q ),
	.prn(vcc));
defparam \out_cnt[0] .is_wysiwyg = "true";
defparam \out_cnt[0] .power_up = "low";

cycloneiv_lcell_comb \out_cnt[3]~0 (
	.dataa(\out_cnt[0]~q ),
	.datab(\out_cnt[1]~q ),
	.datac(\out_cnt[2]~q ),
	.datad(\out_cnt[3]~q ),
	.cin(gnd),
	.combout(\out_cnt[3]~0_combout ),
	.cout());
defparam \out_cnt[3]~0 .lut_mask = 16'h7FFF;
defparam \out_cnt[3]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~1 (
	.dataa(\Equal2~0_combout ),
	.datab(\Equal2~1_combout ),
	.datac(\in_cnt[0]~q ),
	.datad(\gen_out_cnt_p~0_combout ),
	.cin(gnd),
	.combout(\out_cnt[3]~1_combout ),
	.cout());
defparam \out_cnt[3]~1 .lut_mask = 16'h7FFF;
defparam \out_cnt[3]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[3]~2 (
	.dataa(enable),
	.datab(\out_cnt[3]~0_combout ),
	.datac(\out_cnt[3]~1_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_cnt[3]~2_combout ),
	.cout());
defparam \out_cnt[3]~2 .lut_mask = 16'hFDFD;
defparam \out_cnt[3]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_cnt[1]~4 (
	.dataa(\out_cnt[1]~q ),
	.datab(\out_cnt[3]~2_combout ),
	.datac(\out_cnt[3]~3_combout ),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\out_cnt[1]~4_combout ),
	.cout());
defparam \out_cnt[1]~4 .lut_mask = 16'h9F6F;
defparam \out_cnt[1]~4 .sum_lutc_input = "datac";

dffeas \out_cnt[1] (
	.clk(clk),
	.d(\out_cnt[1]~4_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.q(\out_cnt[1]~q ),
	.prn(vcc));
defparam \out_cnt[1] .is_wysiwyg = "true";
defparam \out_cnt[1] .power_up = "low";

cycloneiv_lcell_comb \Equal2~0 (
	.dataa(fftpts_less_one_0),
	.datab(fftpts_less_one_1),
	.datac(\out_cnt[1]~q ),
	.datad(\out_cnt[0]~q ),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
defparam \Equal2~0 .lut_mask = 16'h6996;
defparam \Equal2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \shift~0 (
	.dataa(\gen_out_cnt_p~1_combout ),
	.datab(\shift~q ),
	.datac(\Equal2~0_combout ),
	.datad(\Equal2~1_combout ),
	.cin(gnd),
	.combout(\shift~0_combout ),
	.cout());
defparam \shift~0 .lut_mask = 16'hEFFF;
defparam \shift~0 .sum_lutc_input = "datac";

dffeas shift(
	.clk(clk),
	.d(\shift~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\shift~q ),
	.prn(vcc));
defparam shift.is_wysiwyg = "true";
defparam shift.power_up = "low";

cycloneiv_lcell_comb \out_inverse~0 (
	.dataa(out_inverse1),
	.datab(out_inverse_d_8),
	.datac(\gen_out_cnt_p~1_combout ),
	.datad(enable),
	.cin(gnd),
	.combout(\out_inverse~0_combout ),
	.cout());
defparam \out_inverse~0 .lut_mask = 16'hEFFE;
defparam \out_inverse~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_counter_2 (
	out_stall_d,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	control_s_0,
	out_sop_d_8,
	out_valid_d_8,
	counter_p,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	out_stall_d;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
output 	control_s_0;
input 	out_sop_d_8;
input 	out_valid_d_8;
output 	counter_p;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_s~0_combout ;


dffeas \control_s[0] (
	.clk(clk),
	.d(\control_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(counter_p),
	.q(control_s_0),
	.prn(vcc));
defparam \control_s[0] .is_wysiwyg = "true";
defparam \control_s[0] .power_up = "low";

cycloneiv_lcell_comb \counter_p~0 (
	.dataa(out_valid_d_8),
	.datab(out_valid_s),
	.datac(sop),
	.datad(out_stall_d),
	.cin(gnd),
	.combout(counter_p),
	.cout());
defparam \counter_p~0 .lut_mask = 16'hACFF;
defparam \counter_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~0 (
	.dataa(curr_pwr_2_s),
	.datab(out_sop_d_8),
	.datac(gnd),
	.datad(control_s_0),
	.cin(gnd),
	.combout(\control_s~0_combout ),
	.cout());
defparam \control_s~0 .lut_mask = 16'h9966;
defparam \control_s~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_cma (
	stg_imag_next_0,
	stg_real_next_0,
	stg_imag_next_1,
	stg_real_next_1,
	stg_imag_next_2,
	stg_real_next_2,
	stg_imag_next_3,
	stg_real_next_3,
	stg_imag_next_4,
	stg_real_next_4,
	stg_imag_next_5,
	stg_real_next_5,
	stg_imag_next_6,
	stg_real_next_6,
	stg_imag_next_7,
	stg_real_next_7,
	dataout_2,
	dataout_1,
	dataout_0,
	dataout_21,
	dataout_11,
	dataout_01,
	dataout_3,
	dataout_31,
	dataout_4,
	dataout_41,
	dataout_5,
	dataout_51,
	dataout_6,
	dataout_61,
	dataout_7,
	dataout_71,
	dataout_8,
	dataout_81,
	imagtwid_0,
	imagtwid_1,
	imagtwid_2,
	imagtwid_3,
	imagtwid_4,
	imagtwid_5,
	imagtwid_6,
	imagtwid_7,
	out_stall_d,
	stg_valid_next,
	curr_pwr_2_s,
	sop,
	out_valid_s,
	out_enable,
	stg_inverse_next,
	stg_sop_next,
	out_sop_d_8,
	out_valid_d_8,
	out_inverse_d_8,
	realtwid_0,
	realtwid_1,
	realtwid_2,
	realtwid_3,
	realtwid_4,
	realtwid_5,
	realtwid_6,
	realtwid_7,
	control_s_1,
	control_s_2,
	control_s_0,
	stg_control_next_1,
	stg_control_next_2,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	stg_imag_next_0;
input 	stg_real_next_0;
input 	stg_imag_next_1;
input 	stg_real_next_1;
input 	stg_imag_next_2;
input 	stg_real_next_2;
input 	stg_imag_next_3;
input 	stg_real_next_3;
input 	stg_imag_next_4;
input 	stg_real_next_4;
input 	stg_imag_next_5;
input 	stg_real_next_5;
input 	stg_imag_next_6;
input 	stg_real_next_6;
input 	stg_imag_next_7;
input 	stg_real_next_7;
output 	dataout_2;
output 	dataout_1;
output 	dataout_0;
output 	dataout_21;
output 	dataout_11;
output 	dataout_01;
output 	dataout_3;
output 	dataout_31;
output 	dataout_4;
output 	dataout_41;
output 	dataout_5;
output 	dataout_51;
output 	dataout_6;
output 	dataout_61;
output 	dataout_7;
output 	dataout_71;
output 	dataout_8;
output 	dataout_81;
input 	imagtwid_0;
input 	imagtwid_1;
input 	imagtwid_2;
input 	imagtwid_3;
input 	imagtwid_4;
input 	imagtwid_5;
input 	imagtwid_6;
input 	imagtwid_7;
input 	out_stall_d;
input 	stg_valid_next;
input 	curr_pwr_2_s;
input 	sop;
input 	out_valid_s;
input 	out_enable;
input 	stg_inverse_next;
input 	stg_sop_next;
output 	out_sop_d_8;
output 	out_valid_d_8;
output 	out_inverse_d_8;
input 	realtwid_0;
input 	realtwid_1;
input 	realtwid_2;
input 	realtwid_3;
input 	realtwid_4;
input 	realtwid_5;
input 	realtwid_6;
input 	realtwid_7;
output 	control_s_1;
output 	control_s_2;
output 	control_s_0;
input 	stg_control_next_1;
input 	stg_control_next_2;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:round_imag|conv_round_3:OR_accu~0_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[9]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[8]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[9]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[8]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[10]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[10]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[11]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[11]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[12]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[12]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[13]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[13]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[14]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[14]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:imag_result[15]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:real_result[15]~q ;
wire \imag_result~0_combout ;
wire \imag_result~1_combout ;
wire \imag_result~2_combout ;
wire \imag_result~3_combout ;
wire \imag_result~4_combout ;
wire \imag_result~5_combout ;
wire \imag_result~6_combout ;
wire \imag_result~7_combout ;
wire \imag_result~8_combout ;
wire \imag_result~9_combout ;
wire \real_result~0_combout ;
wire \real_result~1_combout ;
wire \real_result~2_combout ;
wire \real_result~3_combout ;
wire \real_result~4_combout ;
wire \real_result~5_combout ;
wire \real_result~6_combout ;
wire \real_result~7_combout ;
wire \real_result~8_combout ;
wire \real_result~9_combout ;
wire \imag_result~10_combout ;
wire \real_result~10_combout ;
wire \imag_result~11_combout ;
wire \real_result~11_combout ;
wire \imag_result~12_combout ;
wire \real_result~12_combout ;
wire \imag_result~13_combout ;
wire \real_result~13_combout ;
wire \imag_result~14_combout ;
wire \real_result~14_combout ;
wire \imag_result~15_combout ;
wire \real_result~15_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7]~q ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0]~q ;
wire \in_imag_d~0_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1]~q ;
wire \in_imag_d~1_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2]~q ;
wire \in_imag_d~2_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3]~q ;
wire \in_imag_d~3_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4]~q ;
wire \in_imag_d~4_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5]~q ;
wire \in_imag_d~5_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6]~q ;
wire \in_imag_d~6_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7]~q ;
wire \in_imag_d~7_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0]~q ;
wire \in_real_d~0_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1]~q ;
wire \in_real_d~1_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2]~q ;
wire \in_real_d~2_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3]~q ;
wire \in_real_d~3_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4]~q ;
wire \in_real_d~4_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5]~q ;
wire \in_real_d~5_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6]~q ;
wire \in_real_d~6_combout ;
wire \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7]~q ;
wire \in_real_d~7_combout ;
wire \in_imag_dd~0_combout ;
wire \in_imag_dd~1_combout ;
wire \in_imag_dd~2_combout ;
wire \in_imag_dd~3_combout ;
wire \in_imag_dd~4_combout ;
wire \in_imag_dd~5_combout ;
wire \in_imag_dd~6_combout ;
wire \in_imag_dd~7_combout ;
wire \in_real_dd~0_combout ;
wire \in_real_dd~1_combout ;
wire \in_real_dd~2_combout ;
wire \in_real_dd~3_combout ;
wire \in_real_dd~4_combout ;
wire \in_real_dd~5_combout ;
wire \in_real_dd~6_combout ;
wire \in_real_dd~7_combout ;
wire \out_sop_d~9_combout ;
wire \out_sop_d[2]~1_combout ;
wire \out_sop_d[0]~q ;
wire \out_sop_d~8_combout ;
wire \out_sop_d[1]~q ;
wire \out_sop_d~7_combout ;
wire \out_sop_d[2]~q ;
wire \out_sop_d~6_combout ;
wire \out_sop_d[3]~q ;
wire \out_sop_d~5_combout ;
wire \out_sop_d[4]~q ;
wire \out_sop_d~4_combout ;
wire \out_sop_d[5]~q ;
wire \out_sop_d~3_combout ;
wire \out_sop_d[6]~q ;
wire \out_sop_d~2_combout ;
wire \out_sop_d[7]~q ;
wire \out_sop_d~0_combout ;
wire \out_valid_d~8_combout ;
wire \out_valid_d[0]~q ;
wire \out_valid_d~7_combout ;
wire \out_valid_d[1]~q ;
wire \out_valid_d~6_combout ;
wire \out_valid_d[2]~q ;
wire \out_valid_d~5_combout ;
wire \out_valid_d[3]~q ;
wire \out_valid_d~4_combout ;
wire \out_valid_d[4]~q ;
wire \out_valid_d~3_combout ;
wire \out_valid_d[5]~q ;
wire \out_valid_d~2_combout ;
wire \out_valid_d[6]~q ;
wire \out_valid_d~1_combout ;
wire \out_valid_d[7]~q ;
wire \out_valid_d~0_combout ;
wire \out_inverse_d~8_combout ;
wire \out_inverse_d[0]~q ;
wire \out_inverse_d~7_combout ;
wire \out_inverse_d[1]~q ;
wire \out_inverse_d~6_combout ;
wire \out_inverse_d[2]~q ;
wire \out_inverse_d~5_combout ;
wire \out_inverse_d[3]~q ;
wire \out_inverse_d~4_combout ;
wire \out_inverse_d[4]~q ;
wire \out_inverse_d~3_combout ;
wire \out_inverse_d[5]~q ;
wire \out_inverse_d~2_combout ;
wire \out_inverse_d[6]~q ;
wire \out_inverse_d~1_combout ;
wire \out_inverse_d[7]~q ;
wire \out_inverse_d~0_combout ;


ifft_8p_auk_dspip_roundsat \NONA10_C_Mult_Archs:gen_small_mult:round_imag (
	.dataout_2(dataout_2),
	.dataout_1(dataout_1),
	.dataout_0(dataout_0),
	.dataout_3(dataout_3),
	.dataout_4(dataout_4),
	.dataout_5(dataout_5),
	.dataout_6(dataout_6),
	.dataout_7(dataout_7),
	.dataout_8(dataout_8),
	.out_stall_d(out_stall_d),
	.sop(sop),
	.out_valid_s(out_valid_s),
	.out_sop_d_2(\out_sop_d[2]~1_combout ),
	.conv_round_3OR_accu(\NONA10_C_Mult_Archs:gen_small_mult:round_imag|conv_round_3:OR_accu~0_combout ),
	.NONA10_C_Mult_Archsgen_small_multimag_result9(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[9]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result8(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[8]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result7(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[7]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result6(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result3(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result4(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result5(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result0(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result1(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result2(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result10(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[10]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result11(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[11]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result12(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[12]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result13(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[13]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result14(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[14]~q ),
	.NONA10_C_Mult_Archsgen_small_multimag_result15(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[15]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_roundsat_1 \NONA10_C_Mult_Archs:gen_small_mult:round_real (
	.dataout_2(dataout_21),
	.dataout_1(dataout_11),
	.dataout_0(dataout_01),
	.dataout_3(dataout_31),
	.dataout_4(dataout_41),
	.dataout_5(dataout_51),
	.dataout_6(dataout_61),
	.dataout_7(dataout_71),
	.dataout_8(dataout_81),
	.out_sop_d_2(\out_sop_d[2]~1_combout ),
	.reset(\NONA10_C_Mult_Archs:gen_small_mult:round_imag|conv_round_3:OR_accu~0_combout ),
	.NONA10_C_Mult_Archsgen_small_multreal_result9(\NONA10_C_Mult_Archs:gen_small_mult:real_result[9]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result8(\NONA10_C_Mult_Archs:gen_small_mult:real_result[8]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result7(\NONA10_C_Mult_Archs:gen_small_mult:real_result[7]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result6(\NONA10_C_Mult_Archs:gen_small_mult:real_result[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result3(\NONA10_C_Mult_Archs:gen_small_mult:real_result[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result4(\NONA10_C_Mult_Archs:gen_small_mult:real_result[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result5(\NONA10_C_Mult_Archs:gen_small_mult:real_result[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result0(\NONA10_C_Mult_Archs:gen_small_mult:real_result[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result1(\NONA10_C_Mult_Archs:gen_small_mult:real_result[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result2(\NONA10_C_Mult_Archs:gen_small_mult:real_result[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result10(\NONA10_C_Mult_Archs:gen_small_mult:real_result[10]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result11(\NONA10_C_Mult_Archs:gen_small_mult:real_result[11]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result12(\NONA10_C_Mult_Archs:gen_small_mult:real_result[12]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result13(\NONA10_C_Mult_Archs:gen_small_mult:real_result[13]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result14(\NONA10_C_Mult_Archs:gen_small_mult:real_result[14]~q ),
	.NONA10_C_Mult_Archsgen_small_multreal_result15(\NONA10_C_Mult_Archs:gen_small_mult:real_result[15]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_altera_fft_mult_add \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag (
	.dffe5a_9(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.dffe5a_8(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.dffe5a_7(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.dffe5a_6(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.dffe5a_3(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.dffe5a_4(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.dffe5a_5(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.dffe5a_0(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.dffe5a_1(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.dffe5a_2(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.dffe5a_10(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.dffe5a_11(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.dffe5a_12(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.dffe5a_13(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.dffe5a_14(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.dffe5a_15(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.imagtwid_0(imagtwid_0),
	.imagtwid_1(imagtwid_1),
	.imagtwid_2(imagtwid_2),
	.imagtwid_3(imagtwid_3),
	.imagtwid_4(imagtwid_4),
	.imagtwid_5(imagtwid_5),
	.imagtwid_6(imagtwid_6),
	.imagtwid_7(imagtwid_7),
	.out_enable(out_enable),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d0(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d1(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d2(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d3(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d4(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d5(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d6(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d7(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7]~q ),
	.realtwid_0(realtwid_0),
	.realtwid_1(realtwid_1),
	.realtwid_2(realtwid_2),
	.realtwid_3(realtwid_3),
	.realtwid_4(realtwid_4),
	.realtwid_5(realtwid_5),
	.realtwid_6(realtwid_6),
	.realtwid_7(realtwid_7),
	.NONA10_C_Mult_Archsgen_small_multin_real_d0(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d1(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d2(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d3(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d4(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d5(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d6(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d7(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_altera_fft_mult_add_1 \NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real (
	.dffe7a_9(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.dffe7a_8(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.dffe7a_7(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.dffe7a_6(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.dffe7a_3(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.dffe7a_4(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.dffe7a_5(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.dffe7a_0(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.dffe7a_1(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.dffe7a_2(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.dffe7a_10(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.dffe7a_11(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.dffe7a_12(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.dffe7a_13(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.dffe7a_14(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.dffe7a_15(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.imagtwid_0(imagtwid_0),
	.imagtwid_1(imagtwid_1),
	.imagtwid_2(imagtwid_2),
	.imagtwid_3(imagtwid_3),
	.imagtwid_4(imagtwid_4),
	.imagtwid_5(imagtwid_5),
	.imagtwid_6(imagtwid_6),
	.imagtwid_7(imagtwid_7),
	.out_enable(out_enable),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d0(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d1(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d2(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d3(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d4(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d5(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d6(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_imag_d7(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7]~q ),
	.realtwid_0(realtwid_0),
	.realtwid_1(realtwid_1),
	.realtwid_2(realtwid_2),
	.realtwid_3(realtwid_3),
	.realtwid_4(realtwid_4),
	.realtwid_5(realtwid_5),
	.realtwid_6(realtwid_6),
	.realtwid_7(realtwid_7),
	.NONA10_C_Mult_Archsgen_small_multin_real_d0(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d1(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d2(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d3(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d4(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d5(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d6(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6]~q ),
	.NONA10_C_Mult_Archsgen_small_multin_real_d7(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7]~q ),
	.clk(clk),
	.reset_n(reset));

ifft_8p_auk_dspip_r22sdf_counter_3 bf_counter_inst(
	.stg_valid_next(stg_valid_next),
	.curr_pwr_2_s(curr_pwr_2_s),
	.out_enable(out_enable),
	.stg_sop_next(stg_sop_next),
	.control_s_1(control_s_1),
	.control_s_2(control_s_2),
	.control_s_0(control_s_0),
	.stg_control_next_1(stg_control_next_1),
	.stg_control_next_2(stg_control_next_2),
	.clk(clk),
	.reset(reset));

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[9] (
	.clk(clk),
	.d(\imag_result~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[9]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[9] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[9] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[8] (
	.clk(clk),
	.d(\imag_result~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[8]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[8] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[8] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[7] (
	.clk(clk),
	.d(\imag_result~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[7] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[6] (
	.clk(clk),
	.d(\imag_result~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[6] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[3] (
	.clk(clk),
	.d(\imag_result~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[3] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[4] (
	.clk(clk),
	.d(\imag_result~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[4] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[5] (
	.clk(clk),
	.d(\imag_result~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[5] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[0] (
	.clk(clk),
	.d(\imag_result~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[0] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[1] (
	.clk(clk),
	.d(\imag_result~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[1] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[2] (
	.clk(clk),
	.d(\imag_result~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[2] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[9] (
	.clk(clk),
	.d(\real_result~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[9]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[9] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[9] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[8] (
	.clk(clk),
	.d(\real_result~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[8]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[8] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[8] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[7] (
	.clk(clk),
	.d(\real_result~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[7] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[6] (
	.clk(clk),
	.d(\real_result~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[6] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[3] (
	.clk(clk),
	.d(\real_result~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[3] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[4] (
	.clk(clk),
	.d(\real_result~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[4] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[5] (
	.clk(clk),
	.d(\real_result~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[5] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[0] (
	.clk(clk),
	.d(\real_result~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[0] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[1] (
	.clk(clk),
	.d(\real_result~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[1] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[2] (
	.clk(clk),
	.d(\real_result~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[2] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[10] (
	.clk(clk),
	.d(\imag_result~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[10]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[10] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[10] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[10] (
	.clk(clk),
	.d(\real_result~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[10]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[10] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[10] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[11] (
	.clk(clk),
	.d(\imag_result~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[11]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[11] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[11] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[11] (
	.clk(clk),
	.d(\real_result~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[11]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[11] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[11] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[12] (
	.clk(clk),
	.d(\imag_result~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[12]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[12] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[12] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[12] (
	.clk(clk),
	.d(\real_result~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[12]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[12] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[12] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[13] (
	.clk(clk),
	.d(\imag_result~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[13]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[13] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[13] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[13] (
	.clk(clk),
	.d(\real_result~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[13]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[13] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[13] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[14] (
	.clk(clk),
	.d(\imag_result~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[14]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[14] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[14] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[14] (
	.clk(clk),
	.d(\real_result~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[14]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[14] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[14] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:imag_result[15] (
	.clk(clk),
	.d(\imag_result~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:imag_result[15]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[15] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:imag_result[15] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:real_result[15] (
	.clk(clk),
	.d(\real_result~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:real_result[15]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[15] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:real_result[15] .power_up = "low";

cycloneiv_lcell_comb \imag_result~0 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~0_combout ),
	.cout());
defparam \imag_result~0 .lut_mask = 16'hEEEE;
defparam \imag_result~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~1 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~1_combout ),
	.cout());
defparam \imag_result~1 .lut_mask = 16'hEEEE;
defparam \imag_result~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~2 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~2_combout ),
	.cout());
defparam \imag_result~2 .lut_mask = 16'hEEEE;
defparam \imag_result~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~3 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~3_combout ),
	.cout());
defparam \imag_result~3 .lut_mask = 16'hEEEE;
defparam \imag_result~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~4 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~4_combout ),
	.cout());
defparam \imag_result~4 .lut_mask = 16'hEEEE;
defparam \imag_result~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~5 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~5_combout ),
	.cout());
defparam \imag_result~5 .lut_mask = 16'hEEEE;
defparam \imag_result~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~6 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~6_combout ),
	.cout());
defparam \imag_result~6 .lut_mask = 16'hEEEE;
defparam \imag_result~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~7 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~7_combout ),
	.cout());
defparam \imag_result~7 .lut_mask = 16'hEEEE;
defparam \imag_result~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~8 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~8_combout ),
	.cout());
defparam \imag_result~8 .lut_mask = 16'hEEEE;
defparam \imag_result~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~9 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~9_combout ),
	.cout());
defparam \imag_result~9 .lut_mask = 16'hEEEE;
defparam \imag_result~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~0 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[9]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~0_combout ),
	.cout());
defparam \real_result~0 .lut_mask = 16'hEEEE;
defparam \real_result~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~1 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[8]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~1_combout ),
	.cout());
defparam \real_result~1 .lut_mask = 16'hEEEE;
defparam \real_result~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~2 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~2_combout ),
	.cout());
defparam \real_result~2 .lut_mask = 16'hEEEE;
defparam \real_result~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~3 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~3_combout ),
	.cout());
defparam \real_result~3 .lut_mask = 16'hEEEE;
defparam \real_result~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~4 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~4_combout ),
	.cout());
defparam \real_result~4 .lut_mask = 16'hEEEE;
defparam \real_result~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~5 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~5_combout ),
	.cout());
defparam \real_result~5 .lut_mask = 16'hEEEE;
defparam \real_result~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~6 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~6_combout ),
	.cout());
defparam \real_result~6 .lut_mask = 16'hEEEE;
defparam \real_result~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~7 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~7_combout ),
	.cout());
defparam \real_result~7 .lut_mask = 16'hEEEE;
defparam \real_result~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~8 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~8_combout ),
	.cout());
defparam \real_result~8 .lut_mask = 16'hEEEE;
defparam \real_result~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~9 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~9_combout ),
	.cout());
defparam \real_result~9 .lut_mask = 16'hEEEE;
defparam \real_result~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~10 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~10_combout ),
	.cout());
defparam \imag_result~10 .lut_mask = 16'hEEEE;
defparam \imag_result~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~10 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[10]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~10_combout ),
	.cout());
defparam \real_result~10 .lut_mask = 16'hEEEE;
defparam \real_result~10 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~11 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~11_combout ),
	.cout());
defparam \imag_result~11 .lut_mask = 16'hEEEE;
defparam \imag_result~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~11 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[11]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~11_combout ),
	.cout());
defparam \real_result~11 .lut_mask = 16'hEEEE;
defparam \real_result~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~12 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~12_combout ),
	.cout());
defparam \imag_result~12 .lut_mask = 16'hEEEE;
defparam \imag_result~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~12 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[12]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~12_combout ),
	.cout());
defparam \real_result~12 .lut_mask = 16'hEEEE;
defparam \real_result~12 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~13 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~13_combout ),
	.cout());
defparam \imag_result~13 .lut_mask = 16'hEEEE;
defparam \imag_result~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~13 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[13]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~13_combout ),
	.cout());
defparam \real_result~13 .lut_mask = 16'hEEEE;
defparam \real_result~13 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~14 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~14_combout ),
	.cout());
defparam \imag_result~14 .lut_mask = 16'hEEEE;
defparam \imag_result~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~14 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[14]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~14_combout ),
	.cout());
defparam \real_result~14 .lut_mask = 16'hEEEE;
defparam \real_result~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \imag_result~15 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_imag|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe5a[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\imag_result~15_combout ),
	.cout());
defparam \imag_result~15 .lut_mask = 16'hEEEE;
defparam \imag_result~15 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \real_result~15 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:MULT_ADD_real|use_old_mult_add_gen:ALTMULT_ADD_component|ALTMULT_ADD_component|auto_generated|dffe7a[15]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\real_result~15_combout ),
	.cout());
defparam \real_result~15 .lut_mask = 16'hEEEE;
defparam \real_result~15 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0] (
	.clk(clk),
	.d(\in_imag_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[0] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1] (
	.clk(clk),
	.d(\in_imag_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[1] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2] (
	.clk(clk),
	.d(\in_imag_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[2] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3] (
	.clk(clk),
	.d(\in_imag_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[3] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4] (
	.clk(clk),
	.d(\in_imag_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[4] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5] (
	.clk(clk),
	.d(\in_imag_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[5] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6] (
	.clk(clk),
	.d(\in_imag_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[6] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7] (
	.clk(clk),
	.d(\in_imag_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_d[7] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0] (
	.clk(clk),
	.d(\in_real_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[0] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1] (
	.clk(clk),
	.d(\in_real_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[1] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2] (
	.clk(clk),
	.d(\in_real_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[2] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3] (
	.clk(clk),
	.d(\in_real_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[3] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4] (
	.clk(clk),
	.d(\in_real_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[4] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5] (
	.clk(clk),
	.d(\in_real_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[5] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6] (
	.clk(clk),
	.d(\in_real_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[6] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7] (
	.clk(clk),
	.d(\in_real_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_d[7] .power_up = "low";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0] (
	.clk(clk),
	.d(\in_imag_dd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~0 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~0_combout ),
	.cout());
defparam \in_imag_d~0 .lut_mask = 16'hEEEE;
defparam \in_imag_d~0 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1] (
	.clk(clk),
	.d(\in_imag_dd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~1 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~1_combout ),
	.cout());
defparam \in_imag_d~1 .lut_mask = 16'hEEEE;
defparam \in_imag_d~1 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2] (
	.clk(clk),
	.d(\in_imag_dd~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~2 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~2_combout ),
	.cout());
defparam \in_imag_d~2 .lut_mask = 16'hEEEE;
defparam \in_imag_d~2 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3] (
	.clk(clk),
	.d(\in_imag_dd~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~3 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~3_combout ),
	.cout());
defparam \in_imag_d~3 .lut_mask = 16'hEEEE;
defparam \in_imag_d~3 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4] (
	.clk(clk),
	.d(\in_imag_dd~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~4 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~4_combout ),
	.cout());
defparam \in_imag_d~4 .lut_mask = 16'hEEEE;
defparam \in_imag_d~4 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5] (
	.clk(clk),
	.d(\in_imag_dd~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~5 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~5_combout ),
	.cout());
defparam \in_imag_d~5 .lut_mask = 16'hEEEE;
defparam \in_imag_d~5 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6] (
	.clk(clk),
	.d(\in_imag_dd~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~6 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~6_combout ),
	.cout());
defparam \in_imag_d~6 .lut_mask = 16'hEEEE;
defparam \in_imag_d~6 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7] (
	.clk(clk),
	.d(\in_imag_dd~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7] .power_up = "low";

cycloneiv_lcell_comb \in_imag_d~7 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_imag_dd[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_d~7_combout ),
	.cout());
defparam \in_imag_d~7 .lut_mask = 16'hEEEE;
defparam \in_imag_d~7 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0] (
	.clk(clk),
	.d(\in_real_dd~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~0 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~0_combout ),
	.cout());
defparam \in_real_d~0 .lut_mask = 16'hEEEE;
defparam \in_real_d~0 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1] (
	.clk(clk),
	.d(\in_real_dd~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~1 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~1_combout ),
	.cout());
defparam \in_real_d~1 .lut_mask = 16'hEEEE;
defparam \in_real_d~1 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2] (
	.clk(clk),
	.d(\in_real_dd~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~2 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~2_combout ),
	.cout());
defparam \in_real_d~2 .lut_mask = 16'hEEEE;
defparam \in_real_d~2 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3] (
	.clk(clk),
	.d(\in_real_dd~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~3 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~3_combout ),
	.cout());
defparam \in_real_d~3 .lut_mask = 16'hEEEE;
defparam \in_real_d~3 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4] (
	.clk(clk),
	.d(\in_real_dd~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~4 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~4_combout ),
	.cout());
defparam \in_real_d~4 .lut_mask = 16'hEEEE;
defparam \in_real_d~4 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5] (
	.clk(clk),
	.d(\in_real_dd~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~5 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~5_combout ),
	.cout());
defparam \in_real_d~5 .lut_mask = 16'hEEEE;
defparam \in_real_d~5 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6] (
	.clk(clk),
	.d(\in_real_dd~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~6 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~6_combout ),
	.cout());
defparam \in_real_d~6 .lut_mask = 16'hEEEE;
defparam \in_real_d~6 .sum_lutc_input = "datac";

dffeas \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7] (
	.clk(clk),
	.d(\in_real_dd~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7]~q ),
	.prn(vcc));
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7] .is_wysiwyg = "true";
defparam \NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7] .power_up = "low";

cycloneiv_lcell_comb \in_real_d~7 (
	.dataa(reset),
	.datab(\NONA10_C_Mult_Archs:gen_small_mult:in_real_dd[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_d~7_combout ),
	.cout());
defparam \in_real_d~7 .lut_mask = 16'hEEEE;
defparam \in_real_d~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~0 (
	.dataa(reset),
	.datab(stg_imag_next_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~0_combout ),
	.cout());
defparam \in_imag_dd~0 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~1 (
	.dataa(reset),
	.datab(stg_imag_next_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~1_combout ),
	.cout());
defparam \in_imag_dd~1 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~2 (
	.dataa(reset),
	.datab(stg_imag_next_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~2_combout ),
	.cout());
defparam \in_imag_dd~2 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~3 (
	.dataa(reset),
	.datab(stg_imag_next_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~3_combout ),
	.cout());
defparam \in_imag_dd~3 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~4 (
	.dataa(reset),
	.datab(stg_imag_next_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~4_combout ),
	.cout());
defparam \in_imag_dd~4 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~5 (
	.dataa(reset),
	.datab(stg_imag_next_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~5_combout ),
	.cout());
defparam \in_imag_dd~5 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~6 (
	.dataa(reset),
	.datab(stg_imag_next_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~6_combout ),
	.cout());
defparam \in_imag_dd~6 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_imag_dd~7 (
	.dataa(reset),
	.datab(stg_imag_next_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_imag_dd~7_combout ),
	.cout());
defparam \in_imag_dd~7 .lut_mask = 16'hEEEE;
defparam \in_imag_dd~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~0 (
	.dataa(reset),
	.datab(stg_real_next_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~0_combout ),
	.cout());
defparam \in_real_dd~0 .lut_mask = 16'hEEEE;
defparam \in_real_dd~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~1 (
	.dataa(reset),
	.datab(stg_real_next_1),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~1_combout ),
	.cout());
defparam \in_real_dd~1 .lut_mask = 16'hEEEE;
defparam \in_real_dd~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~2 (
	.dataa(reset),
	.datab(stg_real_next_2),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~2_combout ),
	.cout());
defparam \in_real_dd~2 .lut_mask = 16'hEEEE;
defparam \in_real_dd~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~3 (
	.dataa(reset),
	.datab(stg_real_next_3),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~3_combout ),
	.cout());
defparam \in_real_dd~3 .lut_mask = 16'hEEEE;
defparam \in_real_dd~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~4 (
	.dataa(reset),
	.datab(stg_real_next_4),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~4_combout ),
	.cout());
defparam \in_real_dd~4 .lut_mask = 16'hEEEE;
defparam \in_real_dd~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~5 (
	.dataa(reset),
	.datab(stg_real_next_5),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~5_combout ),
	.cout());
defparam \in_real_dd~5 .lut_mask = 16'hEEEE;
defparam \in_real_dd~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~6 (
	.dataa(reset),
	.datab(stg_real_next_6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~6_combout ),
	.cout());
defparam \in_real_dd~6 .lut_mask = 16'hEEEE;
defparam \in_real_dd~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \in_real_dd~7 (
	.dataa(reset),
	.datab(stg_real_next_7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\in_real_dd~7_combout ),
	.cout());
defparam \in_real_dd~7 .lut_mask = 16'hEEEE;
defparam \in_real_dd~7 .sum_lutc_input = "datac";

dffeas \out_sop_d[8] (
	.clk(clk),
	.d(\out_sop_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(out_sop_d_8),
	.prn(vcc));
defparam \out_sop_d[8] .is_wysiwyg = "true";
defparam \out_sop_d[8] .power_up = "low";

dffeas \out_valid_d[8] (
	.clk(clk),
	.d(\out_valid_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(out_valid_d_8),
	.prn(vcc));
defparam \out_valid_d[8] .is_wysiwyg = "true";
defparam \out_valid_d[8] .power_up = "low";

dffeas \out_inverse_d[8] (
	.clk(clk),
	.d(\out_inverse_d~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(out_inverse_d_8),
	.prn(vcc));
defparam \out_inverse_d[8] .is_wysiwyg = "true";
defparam \out_inverse_d[8] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~9 (
	.dataa(reset),
	.datab(stg_sop_next),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~9_combout ),
	.cout());
defparam \out_sop_d~9 .lut_mask = 16'hEEEE;
defparam \out_sop_d~9 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_sop_d[2]~1 (
	.dataa(reset),
	.datab(out_stall_d),
	.datac(sop),
	.datad(out_valid_s),
	.cin(gnd),
	.combout(\out_sop_d[2]~1_combout ),
	.cout());
defparam \out_sop_d[2]~1 .lut_mask = 16'hF737;
defparam \out_sop_d[2]~1 .sum_lutc_input = "datac";

dffeas \out_sop_d[0] (
	.clk(clk),
	.d(\out_sop_d~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[0]~q ),
	.prn(vcc));
defparam \out_sop_d[0] .is_wysiwyg = "true";
defparam \out_sop_d[0] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~8 (
	.dataa(reset),
	.datab(\out_sop_d[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~8_combout ),
	.cout());
defparam \out_sop_d~8 .lut_mask = 16'hEEEE;
defparam \out_sop_d~8 .sum_lutc_input = "datac";

dffeas \out_sop_d[1] (
	.clk(clk),
	.d(\out_sop_d~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[1]~q ),
	.prn(vcc));
defparam \out_sop_d[1] .is_wysiwyg = "true";
defparam \out_sop_d[1] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~7 (
	.dataa(reset),
	.datab(\out_sop_d[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~7_combout ),
	.cout());
defparam \out_sop_d~7 .lut_mask = 16'hEEEE;
defparam \out_sop_d~7 .sum_lutc_input = "datac";

dffeas \out_sop_d[2] (
	.clk(clk),
	.d(\out_sop_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[2]~q ),
	.prn(vcc));
defparam \out_sop_d[2] .is_wysiwyg = "true";
defparam \out_sop_d[2] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~6 (
	.dataa(reset),
	.datab(\out_sop_d[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~6_combout ),
	.cout());
defparam \out_sop_d~6 .lut_mask = 16'hEEEE;
defparam \out_sop_d~6 .sum_lutc_input = "datac";

dffeas \out_sop_d[3] (
	.clk(clk),
	.d(\out_sop_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[3]~q ),
	.prn(vcc));
defparam \out_sop_d[3] .is_wysiwyg = "true";
defparam \out_sop_d[3] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~5 (
	.dataa(reset),
	.datab(\out_sop_d[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~5_combout ),
	.cout());
defparam \out_sop_d~5 .lut_mask = 16'hEEEE;
defparam \out_sop_d~5 .sum_lutc_input = "datac";

dffeas \out_sop_d[4] (
	.clk(clk),
	.d(\out_sop_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[4]~q ),
	.prn(vcc));
defparam \out_sop_d[4] .is_wysiwyg = "true";
defparam \out_sop_d[4] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~4 (
	.dataa(reset),
	.datab(\out_sop_d[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~4_combout ),
	.cout());
defparam \out_sop_d~4 .lut_mask = 16'hEEEE;
defparam \out_sop_d~4 .sum_lutc_input = "datac";

dffeas \out_sop_d[5] (
	.clk(clk),
	.d(\out_sop_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[5]~q ),
	.prn(vcc));
defparam \out_sop_d[5] .is_wysiwyg = "true";
defparam \out_sop_d[5] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~3 (
	.dataa(reset),
	.datab(\out_sop_d[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~3_combout ),
	.cout());
defparam \out_sop_d~3 .lut_mask = 16'hEEEE;
defparam \out_sop_d~3 .sum_lutc_input = "datac";

dffeas \out_sop_d[6] (
	.clk(clk),
	.d(\out_sop_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[6]~q ),
	.prn(vcc));
defparam \out_sop_d[6] .is_wysiwyg = "true";
defparam \out_sop_d[6] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~2 (
	.dataa(reset),
	.datab(\out_sop_d[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~2_combout ),
	.cout());
defparam \out_sop_d~2 .lut_mask = 16'hEEEE;
defparam \out_sop_d~2 .sum_lutc_input = "datac";

dffeas \out_sop_d[7] (
	.clk(clk),
	.d(\out_sop_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_sop_d[7]~q ),
	.prn(vcc));
defparam \out_sop_d[7] .is_wysiwyg = "true";
defparam \out_sop_d[7] .power_up = "low";

cycloneiv_lcell_comb \out_sop_d~0 (
	.dataa(reset),
	.datab(\out_sop_d[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_sop_d~0_combout ),
	.cout());
defparam \out_sop_d~0 .lut_mask = 16'hEEEE;
defparam \out_sop_d~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_valid_d~8 (
	.dataa(reset),
	.datab(curr_pwr_2_s),
	.datac(stg_valid_next),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~8_combout ),
	.cout());
defparam \out_valid_d~8 .lut_mask = 16'hFEFE;
defparam \out_valid_d~8 .sum_lutc_input = "datac";

dffeas \out_valid_d[0] (
	.clk(clk),
	.d(\out_valid_d~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[0]~q ),
	.prn(vcc));
defparam \out_valid_d[0] .is_wysiwyg = "true";
defparam \out_valid_d[0] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~7 (
	.dataa(reset),
	.datab(\out_valid_d[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~7_combout ),
	.cout());
defparam \out_valid_d~7 .lut_mask = 16'hEEEE;
defparam \out_valid_d~7 .sum_lutc_input = "datac";

dffeas \out_valid_d[1] (
	.clk(clk),
	.d(\out_valid_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[1]~q ),
	.prn(vcc));
defparam \out_valid_d[1] .is_wysiwyg = "true";
defparam \out_valid_d[1] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~6 (
	.dataa(reset),
	.datab(\out_valid_d[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~6_combout ),
	.cout());
defparam \out_valid_d~6 .lut_mask = 16'hEEEE;
defparam \out_valid_d~6 .sum_lutc_input = "datac";

dffeas \out_valid_d[2] (
	.clk(clk),
	.d(\out_valid_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[2]~q ),
	.prn(vcc));
defparam \out_valid_d[2] .is_wysiwyg = "true";
defparam \out_valid_d[2] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~5 (
	.dataa(reset),
	.datab(\out_valid_d[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~5_combout ),
	.cout());
defparam \out_valid_d~5 .lut_mask = 16'hEEEE;
defparam \out_valid_d~5 .sum_lutc_input = "datac";

dffeas \out_valid_d[3] (
	.clk(clk),
	.d(\out_valid_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[3]~q ),
	.prn(vcc));
defparam \out_valid_d[3] .is_wysiwyg = "true";
defparam \out_valid_d[3] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~4 (
	.dataa(reset),
	.datab(\out_valid_d[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~4_combout ),
	.cout());
defparam \out_valid_d~4 .lut_mask = 16'hEEEE;
defparam \out_valid_d~4 .sum_lutc_input = "datac";

dffeas \out_valid_d[4] (
	.clk(clk),
	.d(\out_valid_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[4]~q ),
	.prn(vcc));
defparam \out_valid_d[4] .is_wysiwyg = "true";
defparam \out_valid_d[4] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~3 (
	.dataa(reset),
	.datab(\out_valid_d[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~3_combout ),
	.cout());
defparam \out_valid_d~3 .lut_mask = 16'hEEEE;
defparam \out_valid_d~3 .sum_lutc_input = "datac";

dffeas \out_valid_d[5] (
	.clk(clk),
	.d(\out_valid_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[5]~q ),
	.prn(vcc));
defparam \out_valid_d[5] .is_wysiwyg = "true";
defparam \out_valid_d[5] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~2 (
	.dataa(reset),
	.datab(\out_valid_d[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~2_combout ),
	.cout());
defparam \out_valid_d~2 .lut_mask = 16'hEEEE;
defparam \out_valid_d~2 .sum_lutc_input = "datac";

dffeas \out_valid_d[6] (
	.clk(clk),
	.d(\out_valid_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[6]~q ),
	.prn(vcc));
defparam \out_valid_d[6] .is_wysiwyg = "true";
defparam \out_valid_d[6] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~1 (
	.dataa(reset),
	.datab(\out_valid_d[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~1_combout ),
	.cout());
defparam \out_valid_d~1 .lut_mask = 16'hEEEE;
defparam \out_valid_d~1 .sum_lutc_input = "datac";

dffeas \out_valid_d[7] (
	.clk(clk),
	.d(\out_valid_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_valid_d[7]~q ),
	.prn(vcc));
defparam \out_valid_d[7] .is_wysiwyg = "true";
defparam \out_valid_d[7] .power_up = "low";

cycloneiv_lcell_comb \out_valid_d~0 (
	.dataa(reset),
	.datab(\out_valid_d[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_valid_d~0_combout ),
	.cout());
defparam \out_valid_d~0 .lut_mask = 16'hEEEE;
defparam \out_valid_d~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \out_inverse_d~8 (
	.dataa(reset),
	.datab(stg_inverse_next),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~8_combout ),
	.cout());
defparam \out_inverse_d~8 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~8 .sum_lutc_input = "datac";

dffeas \out_inverse_d[0] (
	.clk(clk),
	.d(\out_inverse_d~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[0]~q ),
	.prn(vcc));
defparam \out_inverse_d[0] .is_wysiwyg = "true";
defparam \out_inverse_d[0] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~7 (
	.dataa(reset),
	.datab(\out_inverse_d[0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~7_combout ),
	.cout());
defparam \out_inverse_d~7 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~7 .sum_lutc_input = "datac";

dffeas \out_inverse_d[1] (
	.clk(clk),
	.d(\out_inverse_d~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[1]~q ),
	.prn(vcc));
defparam \out_inverse_d[1] .is_wysiwyg = "true";
defparam \out_inverse_d[1] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~6 (
	.dataa(reset),
	.datab(\out_inverse_d[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~6_combout ),
	.cout());
defparam \out_inverse_d~6 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~6 .sum_lutc_input = "datac";

dffeas \out_inverse_d[2] (
	.clk(clk),
	.d(\out_inverse_d~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[2]~q ),
	.prn(vcc));
defparam \out_inverse_d[2] .is_wysiwyg = "true";
defparam \out_inverse_d[2] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~5 (
	.dataa(reset),
	.datab(\out_inverse_d[2]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~5_combout ),
	.cout());
defparam \out_inverse_d~5 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~5 .sum_lutc_input = "datac";

dffeas \out_inverse_d[3] (
	.clk(clk),
	.d(\out_inverse_d~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[3]~q ),
	.prn(vcc));
defparam \out_inverse_d[3] .is_wysiwyg = "true";
defparam \out_inverse_d[3] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~4 (
	.dataa(reset),
	.datab(\out_inverse_d[3]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~4_combout ),
	.cout());
defparam \out_inverse_d~4 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~4 .sum_lutc_input = "datac";

dffeas \out_inverse_d[4] (
	.clk(clk),
	.d(\out_inverse_d~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[4]~q ),
	.prn(vcc));
defparam \out_inverse_d[4] .is_wysiwyg = "true";
defparam \out_inverse_d[4] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~3 (
	.dataa(reset),
	.datab(\out_inverse_d[4]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~3_combout ),
	.cout());
defparam \out_inverse_d~3 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~3 .sum_lutc_input = "datac";

dffeas \out_inverse_d[5] (
	.clk(clk),
	.d(\out_inverse_d~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[5]~q ),
	.prn(vcc));
defparam \out_inverse_d[5] .is_wysiwyg = "true";
defparam \out_inverse_d[5] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~2 (
	.dataa(reset),
	.datab(\out_inverse_d[5]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~2_combout ),
	.cout());
defparam \out_inverse_d~2 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~2 .sum_lutc_input = "datac";

dffeas \out_inverse_d[6] (
	.clk(clk),
	.d(\out_inverse_d~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[6]~q ),
	.prn(vcc));
defparam \out_inverse_d[6] .is_wysiwyg = "true";
defparam \out_inverse_d[6] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~1 (
	.dataa(reset),
	.datab(\out_inverse_d[6]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~1_combout ),
	.cout());
defparam \out_inverse_d~1 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~1 .sum_lutc_input = "datac";

dffeas \out_inverse_d[7] (
	.clk(clk),
	.d(\out_inverse_d~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\out_sop_d[2]~1_combout ),
	.q(\out_inverse_d[7]~q ),
	.prn(vcc));
defparam \out_inverse_d[7] .is_wysiwyg = "true";
defparam \out_inverse_d[7] .power_up = "low";

cycloneiv_lcell_comb \out_inverse_d~0 (
	.dataa(reset),
	.datab(\out_inverse_d[7]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\out_inverse_d~0_combout ),
	.cout());
defparam \out_inverse_d~0 .lut_mask = 16'hEEEE;
defparam \out_inverse_d~0 .sum_lutc_input = "datac";

endmodule

module ifft_8p_altera_fft_mult_add (
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_3,
	dffe5a_4,
	dffe5a_5,
	dffe5a_0,
	dffe5a_1,
	dffe5a_2,
	dffe5a_10,
	dffe5a_11,
	dffe5a_12,
	dffe5a_13,
	dffe5a_14,
	dffe5a_15,
	imagtwid_0,
	imagtwid_1,
	imagtwid_2,
	imagtwid_3,
	imagtwid_4,
	imagtwid_5,
	imagtwid_6,
	imagtwid_7,
	out_enable,
	NONA10_C_Mult_Archsgen_small_multin_imag_d0,
	NONA10_C_Mult_Archsgen_small_multin_imag_d1,
	NONA10_C_Mult_Archsgen_small_multin_imag_d2,
	NONA10_C_Mult_Archsgen_small_multin_imag_d3,
	NONA10_C_Mult_Archsgen_small_multin_imag_d4,
	NONA10_C_Mult_Archsgen_small_multin_imag_d5,
	NONA10_C_Mult_Archsgen_small_multin_imag_d6,
	NONA10_C_Mult_Archsgen_small_multin_imag_d7,
	realtwid_0,
	realtwid_1,
	realtwid_2,
	realtwid_3,
	realtwid_4,
	realtwid_5,
	realtwid_6,
	realtwid_7,
	NONA10_C_Mult_Archsgen_small_multin_real_d0,
	NONA10_C_Mult_Archsgen_small_multin_real_d1,
	NONA10_C_Mult_Archsgen_small_multin_real_d2,
	NONA10_C_Mult_Archsgen_small_multin_real_d3,
	NONA10_C_Mult_Archsgen_small_multin_real_d4,
	NONA10_C_Mult_Archsgen_small_multin_real_d5,
	NONA10_C_Mult_Archsgen_small_multin_real_d6,
	NONA10_C_Mult_Archsgen_small_multin_real_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_3;
output 	dffe5a_4;
output 	dffe5a_5;
output 	dffe5a_0;
output 	dffe5a_1;
output 	dffe5a_2;
output 	dffe5a_10;
output 	dffe5a_11;
output 	dffe5a_12;
output 	dffe5a_13;
output 	dffe5a_14;
output 	dffe5a_15;
input 	imagtwid_0;
input 	imagtwid_1;
input 	imagtwid_2;
input 	imagtwid_3;
input 	imagtwid_4;
input 	imagtwid_5;
input 	imagtwid_6;
input 	imagtwid_7;
input 	out_enable;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d0;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d1;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d2;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d3;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d4;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d5;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d6;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d7;
input 	realtwid_0;
input 	realtwid_1;
input 	realtwid_2;
input 	realtwid_3;
input 	realtwid_4;
input 	realtwid_5;
input 	realtwid_6;
input 	realtwid_7;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d0;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d1;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d2;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d3;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d4;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d5;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d6;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altera_fft_mult_add_old \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_3(dffe5a_3),
	.dffe5a_4(dffe5a_4),
	.dffe5a_5(dffe5a_5),
	.dffe5a_0(dffe5a_0),
	.dffe5a_1(dffe5a_1),
	.dffe5a_2(dffe5a_2),
	.dffe5a_10(dffe5a_10),
	.dffe5a_11(dffe5a_11),
	.dffe5a_12(dffe5a_12),
	.dffe5a_13(dffe5a_13),
	.dffe5a_14(dffe5a_14),
	.dffe5a_15(dffe5a_15),
	.datab({realtwid_7,realtwid_6,realtwid_5,realtwid_4,realtwid_3,realtwid_2,realtwid_1,realtwid_0,imagtwid_7,imagtwid_6,imagtwid_5,imagtwid_4,imagtwid_3,imagtwid_2,imagtwid_1,imagtwid_0}),
	.ena0(out_enable),
	.dataa({NONA10_C_Mult_Archsgen_small_multin_imag_d7,NONA10_C_Mult_Archsgen_small_multin_imag_d6,NONA10_C_Mult_Archsgen_small_multin_imag_d5,NONA10_C_Mult_Archsgen_small_multin_imag_d4,NONA10_C_Mult_Archsgen_small_multin_imag_d3,
NONA10_C_Mult_Archsgen_small_multin_imag_d2,NONA10_C_Mult_Archsgen_small_multin_imag_d1,NONA10_C_Mult_Archsgen_small_multin_imag_d0,NONA10_C_Mult_Archsgen_small_multin_real_d7,NONA10_C_Mult_Archsgen_small_multin_real_d6,
NONA10_C_Mult_Archsgen_small_multin_real_d5,NONA10_C_Mult_Archsgen_small_multin_real_d4,NONA10_C_Mult_Archsgen_small_multin_real_d3,NONA10_C_Mult_Archsgen_small_multin_real_d2,NONA10_C_Mult_Archsgen_small_multin_real_d1,
NONA10_C_Mult_Archsgen_small_multin_real_d0}),
	.clock0(clk),
	.aclr0(reset_n));

endmodule

module ifft_8p_altera_fft_mult_add_old (
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_3,
	dffe5a_4,
	dffe5a_5,
	dffe5a_0,
	dffe5a_1,
	dffe5a_2,
	dffe5a_10,
	dffe5a_11,
	dffe5a_12,
	dffe5a_13,
	dffe5a_14,
	dffe5a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_3;
output 	dffe5a_4;
output 	dffe5a_5;
output 	dffe5a_0;
output 	dffe5a_1;
output 	dffe5a_2;
output 	dffe5a_10;
output 	dffe5a_11;
output 	dffe5a_12;
output 	dffe5a_13;
output 	dffe5a_14;
output 	dffe5a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altmult_add_1 ALTMULT_ADD_component(
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_3(dffe5a_3),
	.dffe5a_4(dffe5a_4),
	.dffe5a_5(dffe5a_5),
	.dffe5a_0(dffe5a_0),
	.dffe5a_1(dffe5a_1),
	.dffe5a_2(dffe5a_2),
	.dffe5a_10(dffe5a_10),
	.dffe5a_11(dffe5a_11),
	.dffe5a_12(dffe5a_12),
	.dffe5a_13(dffe5a_13),
	.dffe5a_14(dffe5a_14),
	.dffe5a_15(dffe5a_15),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.ena0(ena0),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_altmult_add_1 (
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_3,
	dffe5a_4,
	dffe5a_5,
	dffe5a_0,
	dffe5a_1,
	dffe5a_2,
	dffe5a_10,
	dffe5a_11,
	dffe5a_12,
	dffe5a_13,
	dffe5a_14,
	dffe5a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_3;
output 	dffe5a_4;
output 	dffe5a_5;
output 	dffe5a_0;
output 	dffe5a_1;
output 	dffe5a_2;
output 	dffe5a_10;
output 	dffe5a_11;
output 	dffe5a_12;
output 	dffe5a_13;
output 	dffe5a_14;
output 	dffe5a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_mult_add_1m6g auto_generated(
	.dffe5a_9(dffe5a_9),
	.dffe5a_8(dffe5a_8),
	.dffe5a_7(dffe5a_7),
	.dffe5a_6(dffe5a_6),
	.dffe5a_3(dffe5a_3),
	.dffe5a_4(dffe5a_4),
	.dffe5a_5(dffe5a_5),
	.dffe5a_0(dffe5a_0),
	.dffe5a_1(dffe5a_1),
	.dffe5a_2(dffe5a_2),
	.dffe5a_10(dffe5a_10),
	.dffe5a_11(dffe5a_11),
	.dffe5a_12(dffe5a_12),
	.dffe5a_13(dffe5a_13),
	.dffe5a_14(dffe5a_14),
	.dffe5a_15(dffe5a_15),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.ena0(ena0),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_mult_add_1m6g (
	dffe5a_9,
	dffe5a_8,
	dffe5a_7,
	dffe5a_6,
	dffe5a_3,
	dffe5a_4,
	dffe5a_5,
	dffe5a_0,
	dffe5a_1,
	dffe5a_2,
	dffe5a_10,
	dffe5a_11,
	dffe5a_12,
	dffe5a_13,
	dffe5a_14,
	dffe5a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe5a_9;
output 	dffe5a_8;
output 	dffe5a_7;
output 	dffe5a_6;
output 	dffe5a_3;
output 	dffe5a_4;
output 	dffe5a_5;
output 	dffe5a_0;
output 	dffe5a_1;
output 	dffe5a_2;
output 	dffe5a_10;
output 	dffe5a_11;
output 	dffe5a_12;
output 	dffe5a_13;
output 	dffe5a_14;
output 	dffe5a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \dffe5a[0]~17 ;
wire \dffe5a[1]~19 ;
wire \dffe5a[2]~21 ;
wire \dffe5a[3]~23 ;
wire \dffe5a[4]~25 ;
wire \dffe5a[5]~27 ;
wire \dffe5a[6]~29 ;
wire \dffe5a[7]~31 ;
wire \dffe5a[8]~33 ;
wire \dffe5a[9]~34_combout ;
wire \dffe5a[8]~32_combout ;
wire \dffe5a[7]~30_combout ;
wire \dffe5a[6]~28_combout ;
wire \dffe5a[3]~22_combout ;
wire \dffe5a[4]~24_combout ;
wire \dffe5a[5]~26_combout ;
wire \dffe5a[0]~16_combout ;
wire \dffe5a[1]~18_combout ;
wire \dffe5a[2]~20_combout ;
wire \dffe5a[9]~35 ;
wire \dffe5a[10]~36_combout ;
wire \dffe5a[10]~37 ;
wire \dffe5a[11]~38_combout ;
wire \dffe5a[11]~39 ;
wire \dffe5a[12]~40_combout ;
wire \dffe5a[12]~41 ;
wire \dffe5a[13]~42_combout ;
wire \dffe5a[13]~43 ;
wire \dffe5a[14]~44_combout ;
wire \dffe5a[14]~45 ;
wire \dffe5a[15]~46_combout ;


ifft_8p_ded_mult_hb91_1 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.ena({gnd,gnd,gnd,ena0}),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8]}),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8]}),
	.clock({gnd,gnd,gnd,clock0}),
	.aclr({gnd,gnd,gnd,aclr0}));

ifft_8p_ded_mult_hb91 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.ena({gnd,gnd,gnd,ena0}),
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock({gnd,gnd,gnd,clock0}),
	.aclr({gnd,gnd,gnd,aclr0}));

dffeas \dffe5a[9] (
	.clk(clock0),
	.d(\dffe5a[9]~34_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_9),
	.prn(vcc));
defparam \dffe5a[9] .is_wysiwyg = "true";
defparam \dffe5a[9] .power_up = "low";

dffeas \dffe5a[8] (
	.clk(clock0),
	.d(\dffe5a[8]~32_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_8),
	.prn(vcc));
defparam \dffe5a[8] .is_wysiwyg = "true";
defparam \dffe5a[8] .power_up = "low";

dffeas \dffe5a[7] (
	.clk(clock0),
	.d(\dffe5a[7]~30_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_7),
	.prn(vcc));
defparam \dffe5a[7] .is_wysiwyg = "true";
defparam \dffe5a[7] .power_up = "low";

dffeas \dffe5a[6] (
	.clk(clock0),
	.d(\dffe5a[6]~28_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_6),
	.prn(vcc));
defparam \dffe5a[6] .is_wysiwyg = "true";
defparam \dffe5a[6] .power_up = "low";

dffeas \dffe5a[3] (
	.clk(clock0),
	.d(\dffe5a[3]~22_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_3),
	.prn(vcc));
defparam \dffe5a[3] .is_wysiwyg = "true";
defparam \dffe5a[3] .power_up = "low";

dffeas \dffe5a[4] (
	.clk(clock0),
	.d(\dffe5a[4]~24_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_4),
	.prn(vcc));
defparam \dffe5a[4] .is_wysiwyg = "true";
defparam \dffe5a[4] .power_up = "low";

dffeas \dffe5a[5] (
	.clk(clock0),
	.d(\dffe5a[5]~26_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_5),
	.prn(vcc));
defparam \dffe5a[5] .is_wysiwyg = "true";
defparam \dffe5a[5] .power_up = "low";

dffeas \dffe5a[0] (
	.clk(clock0),
	.d(\dffe5a[0]~16_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_0),
	.prn(vcc));
defparam \dffe5a[0] .is_wysiwyg = "true";
defparam \dffe5a[0] .power_up = "low";

dffeas \dffe5a[1] (
	.clk(clock0),
	.d(\dffe5a[1]~18_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_1),
	.prn(vcc));
defparam \dffe5a[1] .is_wysiwyg = "true";
defparam \dffe5a[1] .power_up = "low";

dffeas \dffe5a[2] (
	.clk(clock0),
	.d(\dffe5a[2]~20_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_2),
	.prn(vcc));
defparam \dffe5a[2] .is_wysiwyg = "true";
defparam \dffe5a[2] .power_up = "low";

dffeas \dffe5a[10] (
	.clk(clock0),
	.d(\dffe5a[10]~36_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_10),
	.prn(vcc));
defparam \dffe5a[10] .is_wysiwyg = "true";
defparam \dffe5a[10] .power_up = "low";

dffeas \dffe5a[11] (
	.clk(clock0),
	.d(\dffe5a[11]~38_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_11),
	.prn(vcc));
defparam \dffe5a[11] .is_wysiwyg = "true";
defparam \dffe5a[11] .power_up = "low";

dffeas \dffe5a[12] (
	.clk(clock0),
	.d(\dffe5a[12]~40_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_12),
	.prn(vcc));
defparam \dffe5a[12] .is_wysiwyg = "true";
defparam \dffe5a[12] .power_up = "low";

dffeas \dffe5a[13] (
	.clk(clock0),
	.d(\dffe5a[13]~42_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_13),
	.prn(vcc));
defparam \dffe5a[13] .is_wysiwyg = "true";
defparam \dffe5a[13] .power_up = "low";

dffeas \dffe5a[14] (
	.clk(clock0),
	.d(\dffe5a[14]~44_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_14),
	.prn(vcc));
defparam \dffe5a[14] .is_wysiwyg = "true";
defparam \dffe5a[14] .power_up = "low";

dffeas \dffe5a[15] (
	.clk(clock0),
	.d(\dffe5a[15]~46_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe5a_15),
	.prn(vcc));
defparam \dffe5a[15] .is_wysiwyg = "true";
defparam \dffe5a[15] .power_up = "low";

cycloneiv_lcell_comb \dffe5a[0]~16 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe5a[0]~16_combout ),
	.cout(\dffe5a[0]~17 ));
defparam \dffe5a[0]~16 .lut_mask = 16'h66EE;
defparam \dffe5a[0]~16 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \dffe5a[1]~18 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[0]~17 ),
	.combout(\dffe5a[1]~18_combout ),
	.cout(\dffe5a[1]~19 ));
defparam \dffe5a[1]~18 .lut_mask = 16'h967F;
defparam \dffe5a[1]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[2]~20 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[1]~19 ),
	.combout(\dffe5a[2]~20_combout ),
	.cout(\dffe5a[2]~21 ));
defparam \dffe5a[2]~20 .lut_mask = 16'h96EF;
defparam \dffe5a[2]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[3]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[2]~21 ),
	.combout(\dffe5a[3]~22_combout ),
	.cout(\dffe5a[3]~23 ));
defparam \dffe5a[3]~22 .lut_mask = 16'h967F;
defparam \dffe5a[3]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[4]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[3]~23 ),
	.combout(\dffe5a[4]~24_combout ),
	.cout(\dffe5a[4]~25 ));
defparam \dffe5a[4]~24 .lut_mask = 16'h96EF;
defparam \dffe5a[4]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[5]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[4]~25 ),
	.combout(\dffe5a[5]~26_combout ),
	.cout(\dffe5a[5]~27 ));
defparam \dffe5a[5]~26 .lut_mask = 16'h967F;
defparam \dffe5a[5]~26 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[6]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[5]~27 ),
	.combout(\dffe5a[6]~28_combout ),
	.cout(\dffe5a[6]~29 ));
defparam \dffe5a[6]~28 .lut_mask = 16'h96EF;
defparam \dffe5a[6]~28 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[7]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[6]~29 ),
	.combout(\dffe5a[7]~30_combout ),
	.cout(\dffe5a[7]~31 ));
defparam \dffe5a[7]~30 .lut_mask = 16'h967F;
defparam \dffe5a[7]~30 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[8]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[7]~31 ),
	.combout(\dffe5a[8]~32_combout ),
	.cout(\dffe5a[8]~33 ));
defparam \dffe5a[8]~32 .lut_mask = 16'h96EF;
defparam \dffe5a[8]~32 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[9]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[8]~33 ),
	.combout(\dffe5a[9]~34_combout ),
	.cout(\dffe5a[9]~35 ));
defparam \dffe5a[9]~34 .lut_mask = 16'h967F;
defparam \dffe5a[9]~34 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[10]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[9]~35 ),
	.combout(\dffe5a[10]~36_combout ),
	.cout(\dffe5a[10]~37 ));
defparam \dffe5a[10]~36 .lut_mask = 16'h96EF;
defparam \dffe5a[10]~36 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[11]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[10]~37 ),
	.combout(\dffe5a[11]~38_combout ),
	.cout(\dffe5a[11]~39 ));
defparam \dffe5a[11]~38 .lut_mask = 16'h967F;
defparam \dffe5a[11]~38 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[12]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[11]~39 ),
	.combout(\dffe5a[12]~40_combout ),
	.cout(\dffe5a[12]~41 ));
defparam \dffe5a[12]~40 .lut_mask = 16'h96EF;
defparam \dffe5a[12]~40 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[13]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[12]~41 ),
	.combout(\dffe5a[13]~42_combout ),
	.cout(\dffe5a[13]~43 ));
defparam \dffe5a[13]~42 .lut_mask = 16'h967F;
defparam \dffe5a[13]~42 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[14]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe5a[13]~43 ),
	.combout(\dffe5a[14]~44_combout ),
	.cout(\dffe5a[14]~45 ));
defparam \dffe5a[14]~44 .lut_mask = 16'h96EF;
defparam \dffe5a[14]~44 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe5a[15]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe5a[14]~45 ),
	.combout(\dffe5a[15]~46_combout ),
	.cout());
defparam \dffe5a[15]~46 .lut_mask = 16'h9696;
defparam \dffe5a[15]~46 .sum_lutc_input = "cin";

endmodule

module ifft_8p_ded_mult_hb91 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	datab,
	ena,
	dataa,
	clock,
	aclr)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
input 	[7:0] datab;
input 	[3:0] ena;
input 	[7:0] dataa;
input 	[3:0] clock;
input 	[3:0] aclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];

cycloneiv_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,
\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 16;
defparam mac_out9.output_clock = "0";

cycloneiv_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 8;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 8;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module ifft_8p_ded_mult_hb91_1 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	ena,
	dataa,
	datab,
	clock,
	aclr)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
input 	[3:0] ena;
input 	[7:0] dataa;
input 	[7:0] datab;
input 	[3:0] clock;
input 	[3:0] aclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];

cycloneiv_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,
\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 16;
defparam mac_out9.output_clock = "0";

cycloneiv_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 8;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 8;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module ifft_8p_altera_fft_mult_add_1 (
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_3,
	dffe7a_4,
	dffe7a_5,
	dffe7a_0,
	dffe7a_1,
	dffe7a_2,
	dffe7a_10,
	dffe7a_11,
	dffe7a_12,
	dffe7a_13,
	dffe7a_14,
	dffe7a_15,
	imagtwid_0,
	imagtwid_1,
	imagtwid_2,
	imagtwid_3,
	imagtwid_4,
	imagtwid_5,
	imagtwid_6,
	imagtwid_7,
	out_enable,
	NONA10_C_Mult_Archsgen_small_multin_imag_d0,
	NONA10_C_Mult_Archsgen_small_multin_imag_d1,
	NONA10_C_Mult_Archsgen_small_multin_imag_d2,
	NONA10_C_Mult_Archsgen_small_multin_imag_d3,
	NONA10_C_Mult_Archsgen_small_multin_imag_d4,
	NONA10_C_Mult_Archsgen_small_multin_imag_d5,
	NONA10_C_Mult_Archsgen_small_multin_imag_d6,
	NONA10_C_Mult_Archsgen_small_multin_imag_d7,
	realtwid_0,
	realtwid_1,
	realtwid_2,
	realtwid_3,
	realtwid_4,
	realtwid_5,
	realtwid_6,
	realtwid_7,
	NONA10_C_Mult_Archsgen_small_multin_real_d0,
	NONA10_C_Mult_Archsgen_small_multin_real_d1,
	NONA10_C_Mult_Archsgen_small_multin_real_d2,
	NONA10_C_Mult_Archsgen_small_multin_real_d3,
	NONA10_C_Mult_Archsgen_small_multin_real_d4,
	NONA10_C_Mult_Archsgen_small_multin_real_d5,
	NONA10_C_Mult_Archsgen_small_multin_real_d6,
	NONA10_C_Mult_Archsgen_small_multin_real_d7,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_3;
output 	dffe7a_4;
output 	dffe7a_5;
output 	dffe7a_0;
output 	dffe7a_1;
output 	dffe7a_2;
output 	dffe7a_10;
output 	dffe7a_11;
output 	dffe7a_12;
output 	dffe7a_13;
output 	dffe7a_14;
output 	dffe7a_15;
input 	imagtwid_0;
input 	imagtwid_1;
input 	imagtwid_2;
input 	imagtwid_3;
input 	imagtwid_4;
input 	imagtwid_5;
input 	imagtwid_6;
input 	imagtwid_7;
input 	out_enable;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d0;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d1;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d2;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d3;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d4;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d5;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d6;
input 	NONA10_C_Mult_Archsgen_small_multin_imag_d7;
input 	realtwid_0;
input 	realtwid_1;
input 	realtwid_2;
input 	realtwid_3;
input 	realtwid_4;
input 	realtwid_5;
input 	realtwid_6;
input 	realtwid_7;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d0;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d1;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d2;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d3;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d4;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d5;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d6;
input 	NONA10_C_Mult_Archsgen_small_multin_real_d7;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altera_fft_mult_add_old_1 \use_old_mult_add_gen:ALTMULT_ADD_component (
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_3(dffe7a_3),
	.dffe7a_4(dffe7a_4),
	.dffe7a_5(dffe7a_5),
	.dffe7a_0(dffe7a_0),
	.dffe7a_1(dffe7a_1),
	.dffe7a_2(dffe7a_2),
	.dffe7a_10(dffe7a_10),
	.dffe7a_11(dffe7a_11),
	.dffe7a_12(dffe7a_12),
	.dffe7a_13(dffe7a_13),
	.dffe7a_14(dffe7a_14),
	.dffe7a_15(dffe7a_15),
	.datab({imagtwid_7,imagtwid_6,imagtwid_5,imagtwid_4,imagtwid_3,imagtwid_2,imagtwid_1,imagtwid_0,realtwid_7,realtwid_6,realtwid_5,realtwid_4,realtwid_3,realtwid_2,realtwid_1,realtwid_0}),
	.ena0(out_enable),
	.dataa({NONA10_C_Mult_Archsgen_small_multin_imag_d7,NONA10_C_Mult_Archsgen_small_multin_imag_d6,NONA10_C_Mult_Archsgen_small_multin_imag_d5,NONA10_C_Mult_Archsgen_small_multin_imag_d4,NONA10_C_Mult_Archsgen_small_multin_imag_d3,
NONA10_C_Mult_Archsgen_small_multin_imag_d2,NONA10_C_Mult_Archsgen_small_multin_imag_d1,NONA10_C_Mult_Archsgen_small_multin_imag_d0,NONA10_C_Mult_Archsgen_small_multin_real_d7,NONA10_C_Mult_Archsgen_small_multin_real_d6,
NONA10_C_Mult_Archsgen_small_multin_real_d5,NONA10_C_Mult_Archsgen_small_multin_real_d4,NONA10_C_Mult_Archsgen_small_multin_real_d3,NONA10_C_Mult_Archsgen_small_multin_real_d2,NONA10_C_Mult_Archsgen_small_multin_real_d1,
NONA10_C_Mult_Archsgen_small_multin_real_d0}),
	.clock0(clk),
	.aclr0(reset_n));

endmodule

module ifft_8p_altera_fft_mult_add_old_1 (
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_3,
	dffe7a_4,
	dffe7a_5,
	dffe7a_0,
	dffe7a_1,
	dffe7a_2,
	dffe7a_10,
	dffe7a_11,
	dffe7a_12,
	dffe7a_13,
	dffe7a_14,
	dffe7a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_3;
output 	dffe7a_4;
output 	dffe7a_5;
output 	dffe7a_0;
output 	dffe7a_1;
output 	dffe7a_2;
output 	dffe7a_10;
output 	dffe7a_11;
output 	dffe7a_12;
output 	dffe7a_13;
output 	dffe7a_14;
output 	dffe7a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altmult_add_2 ALTMULT_ADD_component(
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_3(dffe7a_3),
	.dffe7a_4(dffe7a_4),
	.dffe7a_5(dffe7a_5),
	.dffe7a_0(dffe7a_0),
	.dffe7a_1(dffe7a_1),
	.dffe7a_2(dffe7a_2),
	.dffe7a_10(dffe7a_10),
	.dffe7a_11(dffe7a_11),
	.dffe7a_12(dffe7a_12),
	.dffe7a_13(dffe7a_13),
	.dffe7a_14(dffe7a_14),
	.dffe7a_15(dffe7a_15),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.ena0(ena0),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_altmult_add_2 (
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_3,
	dffe7a_4,
	dffe7a_5,
	dffe7a_0,
	dffe7a_1,
	dffe7a_2,
	dffe7a_10,
	dffe7a_11,
	dffe7a_12,
	dffe7a_13,
	dffe7a_14,
	dffe7a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_3;
output 	dffe7a_4;
output 	dffe7a_5;
output 	dffe7a_0;
output 	dffe7a_1;
output 	dffe7a_2;
output 	dffe7a_10;
output 	dffe7a_11;
output 	dffe7a_12;
output 	dffe7a_13;
output 	dffe7a_14;
output 	dffe7a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_mult_add_2n6g auto_generated(
	.dffe7a_9(dffe7a_9),
	.dffe7a_8(dffe7a_8),
	.dffe7a_7(dffe7a_7),
	.dffe7a_6(dffe7a_6),
	.dffe7a_3(dffe7a_3),
	.dffe7a_4(dffe7a_4),
	.dffe7a_5(dffe7a_5),
	.dffe7a_0(dffe7a_0),
	.dffe7a_1(dffe7a_1),
	.dffe7a_2(dffe7a_2),
	.dffe7a_10(dffe7a_10),
	.dffe7a_11(dffe7a_11),
	.dffe7a_12(dffe7a_12),
	.dffe7a_13(dffe7a_13),
	.dffe7a_14(dffe7a_14),
	.dffe7a_15(dffe7a_15),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8],datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.ena0(ena0),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8],dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_mult_add_2n6g (
	dffe7a_9,
	dffe7a_8,
	dffe7a_7,
	dffe7a_6,
	dffe7a_3,
	dffe7a_4,
	dffe7a_5,
	dffe7a_0,
	dffe7a_1,
	dffe7a_2,
	dffe7a_10,
	dffe7a_11,
	dffe7a_12,
	dffe7a_13,
	dffe7a_14,
	dffe7a_15,
	datab,
	ena0,
	dataa,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	dffe7a_9;
output 	dffe7a_8;
output 	dffe7a_7;
output 	dffe7a_6;
output 	dffe7a_3;
output 	dffe7a_4;
output 	dffe7a_5;
output 	dffe7a_0;
output 	dffe7a_1;
output 	dffe7a_2;
output 	dffe7a_10;
output 	dffe7a_11;
output 	dffe7a_12;
output 	dffe7a_13;
output 	dffe7a_14;
output 	dffe7a_15;
input 	[15:0] datab;
input 	ena0;
input 	[15:0] dataa;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \ded_mult2|mac_out9~dataout ;
wire \ded_mult2|mac_out9~DATAOUT1 ;
wire \ded_mult2|mac_out9~DATAOUT2 ;
wire \ded_mult2|mac_out9~DATAOUT3 ;
wire \ded_mult2|mac_out9~DATAOUT4 ;
wire \ded_mult2|mac_out9~DATAOUT5 ;
wire \ded_mult2|mac_out9~DATAOUT6 ;
wire \ded_mult2|mac_out9~DATAOUT7 ;
wire \ded_mult2|mac_out9~DATAOUT8 ;
wire \ded_mult2|mac_out9~DATAOUT9 ;
wire \ded_mult2|mac_out9~DATAOUT10 ;
wire \ded_mult2|mac_out9~DATAOUT11 ;
wire \ded_mult2|mac_out9~DATAOUT12 ;
wire \ded_mult2|mac_out9~DATAOUT13 ;
wire \ded_mult2|mac_out9~DATAOUT14 ;
wire \ded_mult2|mac_out9~DATAOUT15 ;
wire \ded_mult1|mac_out9~dataout ;
wire \ded_mult1|mac_out9~DATAOUT1 ;
wire \ded_mult1|mac_out9~DATAOUT2 ;
wire \ded_mult1|mac_out9~DATAOUT3 ;
wire \ded_mult1|mac_out9~DATAOUT4 ;
wire \ded_mult1|mac_out9~DATAOUT5 ;
wire \ded_mult1|mac_out9~DATAOUT6 ;
wire \ded_mult1|mac_out9~DATAOUT7 ;
wire \ded_mult1|mac_out9~DATAOUT8 ;
wire \ded_mult1|mac_out9~DATAOUT9 ;
wire \ded_mult1|mac_out9~DATAOUT10 ;
wire \ded_mult1|mac_out9~DATAOUT11 ;
wire \ded_mult1|mac_out9~DATAOUT12 ;
wire \ded_mult1|mac_out9~DATAOUT13 ;
wire \ded_mult1|mac_out9~DATAOUT14 ;
wire \ded_mult1|mac_out9~DATAOUT15 ;
wire \dffe7a[0]~17 ;
wire \dffe7a[1]~19 ;
wire \dffe7a[2]~21 ;
wire \dffe7a[3]~23 ;
wire \dffe7a[4]~25 ;
wire \dffe7a[5]~27 ;
wire \dffe7a[6]~29 ;
wire \dffe7a[7]~31 ;
wire \dffe7a[8]~33 ;
wire \dffe7a[9]~34_combout ;
wire \dffe7a[8]~32_combout ;
wire \dffe7a[7]~30_combout ;
wire \dffe7a[6]~28_combout ;
wire \dffe7a[3]~22_combout ;
wire \dffe7a[4]~24_combout ;
wire \dffe7a[5]~26_combout ;
wire \dffe7a[0]~16_combout ;
wire \dffe7a[1]~18_combout ;
wire \dffe7a[2]~20_combout ;
wire \dffe7a[9]~35 ;
wire \dffe7a[10]~36_combout ;
wire \dffe7a[10]~37 ;
wire \dffe7a[11]~38_combout ;
wire \dffe7a[11]~39 ;
wire \dffe7a[12]~40_combout ;
wire \dffe7a[12]~41 ;
wire \dffe7a[13]~42_combout ;
wire \dffe7a[13]~43 ;
wire \dffe7a[14]~44_combout ;
wire \dffe7a[14]~45 ;
wire \dffe7a[15]~46_combout ;


ifft_8p_ded_mult_hb91_3 ded_mult2(
	.mac_out91(\ded_mult2|mac_out9~dataout ),
	.mac_out92(\ded_mult2|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult2|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult2|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult2|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult2|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult2|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult2|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult2|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult2|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult2|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult2|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult2|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult2|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult2|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab({datab[15],datab[14],datab[13],datab[12],datab[11],datab[10],datab[9],datab[8]}),
	.ena({gnd,gnd,gnd,ena0}),
	.dataa({dataa[15],dataa[14],dataa[13],dataa[12],dataa[11],dataa[10],dataa[9],dataa[8]}),
	.clock({gnd,gnd,gnd,clock0}),
	.aclr({gnd,gnd,gnd,aclr0}));

ifft_8p_ded_mult_hb91_2 ded_mult1(
	.mac_out91(\ded_mult1|mac_out9~dataout ),
	.mac_out92(\ded_mult1|mac_out9~DATAOUT1 ),
	.mac_out93(\ded_mult1|mac_out9~DATAOUT2 ),
	.mac_out94(\ded_mult1|mac_out9~DATAOUT3 ),
	.mac_out95(\ded_mult1|mac_out9~DATAOUT4 ),
	.mac_out96(\ded_mult1|mac_out9~DATAOUT5 ),
	.mac_out97(\ded_mult1|mac_out9~DATAOUT6 ),
	.mac_out98(\ded_mult1|mac_out9~DATAOUT7 ),
	.mac_out99(\ded_mult1|mac_out9~DATAOUT8 ),
	.mac_out910(\ded_mult1|mac_out9~DATAOUT9 ),
	.mac_out911(\ded_mult1|mac_out9~DATAOUT10 ),
	.mac_out912(\ded_mult1|mac_out9~DATAOUT11 ),
	.mac_out913(\ded_mult1|mac_out9~DATAOUT12 ),
	.mac_out914(\ded_mult1|mac_out9~DATAOUT13 ),
	.mac_out915(\ded_mult1|mac_out9~DATAOUT14 ),
	.mac_out916(\ded_mult1|mac_out9~DATAOUT15 ),
	.ena({gnd,gnd,gnd,ena0}),
	.datab({datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataa({dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.clock({gnd,gnd,gnd,clock0}),
	.aclr({gnd,gnd,gnd,aclr0}));

dffeas \dffe7a[9] (
	.clk(clock0),
	.d(\dffe7a[9]~34_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_9),
	.prn(vcc));
defparam \dffe7a[9] .is_wysiwyg = "true";
defparam \dffe7a[9] .power_up = "low";

dffeas \dffe7a[8] (
	.clk(clock0),
	.d(\dffe7a[8]~32_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_8),
	.prn(vcc));
defparam \dffe7a[8] .is_wysiwyg = "true";
defparam \dffe7a[8] .power_up = "low";

dffeas \dffe7a[7] (
	.clk(clock0),
	.d(\dffe7a[7]~30_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_7),
	.prn(vcc));
defparam \dffe7a[7] .is_wysiwyg = "true";
defparam \dffe7a[7] .power_up = "low";

dffeas \dffe7a[6] (
	.clk(clock0),
	.d(\dffe7a[6]~28_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_6),
	.prn(vcc));
defparam \dffe7a[6] .is_wysiwyg = "true";
defparam \dffe7a[6] .power_up = "low";

dffeas \dffe7a[3] (
	.clk(clock0),
	.d(\dffe7a[3]~22_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_3),
	.prn(vcc));
defparam \dffe7a[3] .is_wysiwyg = "true";
defparam \dffe7a[3] .power_up = "low";

dffeas \dffe7a[4] (
	.clk(clock0),
	.d(\dffe7a[4]~24_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_4),
	.prn(vcc));
defparam \dffe7a[4] .is_wysiwyg = "true";
defparam \dffe7a[4] .power_up = "low";

dffeas \dffe7a[5] (
	.clk(clock0),
	.d(\dffe7a[5]~26_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_5),
	.prn(vcc));
defparam \dffe7a[5] .is_wysiwyg = "true";
defparam \dffe7a[5] .power_up = "low";

dffeas \dffe7a[0] (
	.clk(clock0),
	.d(\dffe7a[0]~16_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_0),
	.prn(vcc));
defparam \dffe7a[0] .is_wysiwyg = "true";
defparam \dffe7a[0] .power_up = "low";

dffeas \dffe7a[1] (
	.clk(clock0),
	.d(\dffe7a[1]~18_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_1),
	.prn(vcc));
defparam \dffe7a[1] .is_wysiwyg = "true";
defparam \dffe7a[1] .power_up = "low";

dffeas \dffe7a[2] (
	.clk(clock0),
	.d(\dffe7a[2]~20_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_2),
	.prn(vcc));
defparam \dffe7a[2] .is_wysiwyg = "true";
defparam \dffe7a[2] .power_up = "low";

dffeas \dffe7a[10] (
	.clk(clock0),
	.d(\dffe7a[10]~36_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_10),
	.prn(vcc));
defparam \dffe7a[10] .is_wysiwyg = "true";
defparam \dffe7a[10] .power_up = "low";

dffeas \dffe7a[11] (
	.clk(clock0),
	.d(\dffe7a[11]~38_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_11),
	.prn(vcc));
defparam \dffe7a[11] .is_wysiwyg = "true";
defparam \dffe7a[11] .power_up = "low";

dffeas \dffe7a[12] (
	.clk(clock0),
	.d(\dffe7a[12]~40_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_12),
	.prn(vcc));
defparam \dffe7a[12] .is_wysiwyg = "true";
defparam \dffe7a[12] .power_up = "low";

dffeas \dffe7a[13] (
	.clk(clock0),
	.d(\dffe7a[13]~42_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_13),
	.prn(vcc));
defparam \dffe7a[13] .is_wysiwyg = "true";
defparam \dffe7a[13] .power_up = "low";

dffeas \dffe7a[14] (
	.clk(clock0),
	.d(\dffe7a[14]~44_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_14),
	.prn(vcc));
defparam \dffe7a[14] .is_wysiwyg = "true";
defparam \dffe7a[14] .power_up = "low";

dffeas \dffe7a[15] (
	.clk(clock0),
	.d(\dffe7a[15]~46_combout ),
	.asdata(vcc),
	.clrn(aclr0),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(ena0),
	.q(dffe7a_15),
	.prn(vcc));
defparam \dffe7a[15] .is_wysiwyg = "true";
defparam \dffe7a[15] .power_up = "low";

cycloneiv_lcell_comb \dffe7a[0]~16 (
	.dataa(\ded_mult2|mac_out9~dataout ),
	.datab(\ded_mult1|mac_out9~dataout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\dffe7a[0]~16_combout ),
	.cout(\dffe7a[0]~17 ));
defparam \dffe7a[0]~16 .lut_mask = 16'h66DD;
defparam \dffe7a[0]~16 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \dffe7a[1]~18 (
	.dataa(\ded_mult2|mac_out9~DATAOUT1 ),
	.datab(\ded_mult1|mac_out9~DATAOUT1 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[0]~17 ),
	.combout(\dffe7a[1]~18_combout ),
	.cout(\dffe7a[1]~19 ));
defparam \dffe7a[1]~18 .lut_mask = 16'h96BF;
defparam \dffe7a[1]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[2]~20 (
	.dataa(\ded_mult2|mac_out9~DATAOUT2 ),
	.datab(\ded_mult1|mac_out9~DATAOUT2 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[1]~19 ),
	.combout(\dffe7a[2]~20_combout ),
	.cout(\dffe7a[2]~21 ));
defparam \dffe7a[2]~20 .lut_mask = 16'h96DF;
defparam \dffe7a[2]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[3]~22 (
	.dataa(\ded_mult2|mac_out9~DATAOUT3 ),
	.datab(\ded_mult1|mac_out9~DATAOUT3 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[2]~21 ),
	.combout(\dffe7a[3]~22_combout ),
	.cout(\dffe7a[3]~23 ));
defparam \dffe7a[3]~22 .lut_mask = 16'h96BF;
defparam \dffe7a[3]~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[4]~24 (
	.dataa(\ded_mult2|mac_out9~DATAOUT4 ),
	.datab(\ded_mult1|mac_out9~DATAOUT4 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[3]~23 ),
	.combout(\dffe7a[4]~24_combout ),
	.cout(\dffe7a[4]~25 ));
defparam \dffe7a[4]~24 .lut_mask = 16'h96DF;
defparam \dffe7a[4]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[5]~26 (
	.dataa(\ded_mult2|mac_out9~DATAOUT5 ),
	.datab(\ded_mult1|mac_out9~DATAOUT5 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[4]~25 ),
	.combout(\dffe7a[5]~26_combout ),
	.cout(\dffe7a[5]~27 ));
defparam \dffe7a[5]~26 .lut_mask = 16'h96BF;
defparam \dffe7a[5]~26 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[6]~28 (
	.dataa(\ded_mult2|mac_out9~DATAOUT6 ),
	.datab(\ded_mult1|mac_out9~DATAOUT6 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[5]~27 ),
	.combout(\dffe7a[6]~28_combout ),
	.cout(\dffe7a[6]~29 ));
defparam \dffe7a[6]~28 .lut_mask = 16'h96DF;
defparam \dffe7a[6]~28 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[7]~30 (
	.dataa(\ded_mult2|mac_out9~DATAOUT7 ),
	.datab(\ded_mult1|mac_out9~DATAOUT7 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[6]~29 ),
	.combout(\dffe7a[7]~30_combout ),
	.cout(\dffe7a[7]~31 ));
defparam \dffe7a[7]~30 .lut_mask = 16'h96BF;
defparam \dffe7a[7]~30 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[8]~32 (
	.dataa(\ded_mult2|mac_out9~DATAOUT8 ),
	.datab(\ded_mult1|mac_out9~DATAOUT8 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[7]~31 ),
	.combout(\dffe7a[8]~32_combout ),
	.cout(\dffe7a[8]~33 ));
defparam \dffe7a[8]~32 .lut_mask = 16'h96DF;
defparam \dffe7a[8]~32 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[9]~34 (
	.dataa(\ded_mult2|mac_out9~DATAOUT9 ),
	.datab(\ded_mult1|mac_out9~DATAOUT9 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[8]~33 ),
	.combout(\dffe7a[9]~34_combout ),
	.cout(\dffe7a[9]~35 ));
defparam \dffe7a[9]~34 .lut_mask = 16'h96BF;
defparam \dffe7a[9]~34 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[10]~36 (
	.dataa(\ded_mult2|mac_out9~DATAOUT10 ),
	.datab(\ded_mult1|mac_out9~DATAOUT10 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[9]~35 ),
	.combout(\dffe7a[10]~36_combout ),
	.cout(\dffe7a[10]~37 ));
defparam \dffe7a[10]~36 .lut_mask = 16'h96DF;
defparam \dffe7a[10]~36 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[11]~38 (
	.dataa(\ded_mult2|mac_out9~DATAOUT11 ),
	.datab(\ded_mult1|mac_out9~DATAOUT11 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[10]~37 ),
	.combout(\dffe7a[11]~38_combout ),
	.cout(\dffe7a[11]~39 ));
defparam \dffe7a[11]~38 .lut_mask = 16'h96BF;
defparam \dffe7a[11]~38 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[12]~40 (
	.dataa(\ded_mult2|mac_out9~DATAOUT12 ),
	.datab(\ded_mult1|mac_out9~DATAOUT12 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[11]~39 ),
	.combout(\dffe7a[12]~40_combout ),
	.cout(\dffe7a[12]~41 ));
defparam \dffe7a[12]~40 .lut_mask = 16'h96DF;
defparam \dffe7a[12]~40 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[13]~42 (
	.dataa(\ded_mult2|mac_out9~DATAOUT13 ),
	.datab(\ded_mult1|mac_out9~DATAOUT13 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[12]~41 ),
	.combout(\dffe7a[13]~42_combout ),
	.cout(\dffe7a[13]~43 ));
defparam \dffe7a[13]~42 .lut_mask = 16'h96BF;
defparam \dffe7a[13]~42 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[14]~44 (
	.dataa(\ded_mult2|mac_out9~DATAOUT14 ),
	.datab(\ded_mult1|mac_out9~DATAOUT14 ),
	.datac(gnd),
	.datad(vcc),
	.cin(\dffe7a[13]~43 ),
	.combout(\dffe7a[14]~44_combout ),
	.cout(\dffe7a[14]~45 ));
defparam \dffe7a[14]~44 .lut_mask = 16'h96DF;
defparam \dffe7a[14]~44 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \dffe7a[15]~46 (
	.dataa(\ded_mult2|mac_out9~DATAOUT15 ),
	.datab(\ded_mult1|mac_out9~DATAOUT15 ),
	.datac(gnd),
	.datad(gnd),
	.cin(\dffe7a[14]~45 ),
	.combout(\dffe7a[15]~46_combout ),
	.cout());
defparam \dffe7a[15]~46 .lut_mask = 16'h9696;
defparam \dffe7a[15]~46 .sum_lutc_input = "cin";

endmodule

module ifft_8p_ded_mult_hb91_2 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	ena,
	datab,
	dataa,
	clock,
	aclr)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
input 	[3:0] ena;
input 	[7:0] datab;
input 	[7:0] dataa;
input 	[3:0] clock;
input 	[3:0] aclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];

cycloneiv_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,
\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 16;
defparam mac_out9.output_clock = "0";

cycloneiv_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 8;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 8;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module ifft_8p_ded_mult_hb91_3 (
	mac_out91,
	mac_out92,
	mac_out93,
	mac_out94,
	mac_out95,
	mac_out96,
	mac_out97,
	mac_out98,
	mac_out99,
	mac_out910,
	mac_out911,
	mac_out912,
	mac_out913,
	mac_out914,
	mac_out915,
	mac_out916,
	datab,
	ena,
	dataa,
	clock,
	aclr)/* synthesis synthesis_greybox=1 */;
output 	mac_out91;
output 	mac_out92;
output 	mac_out93;
output 	mac_out94;
output 	mac_out95;
output 	mac_out96;
output 	mac_out97;
output 	mac_out98;
output 	mac_out99;
output 	mac_out910;
output 	mac_out911;
output 	mac_out912;
output 	mac_out913;
output 	mac_out914;
output 	mac_out915;
output 	mac_out916;
input 	[7:0] datab;
input 	[3:0] ena;
input 	[7:0] dataa;
input 	[3:0] clock;
input 	[3:0] aclr;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \mac_mult8~dataout ;
wire \mac_mult8~DATAOUT1 ;
wire \mac_mult8~DATAOUT2 ;
wire \mac_mult8~DATAOUT3 ;
wire \mac_mult8~DATAOUT4 ;
wire \mac_mult8~DATAOUT5 ;
wire \mac_mult8~DATAOUT6 ;
wire \mac_mult8~DATAOUT7 ;
wire \mac_mult8~DATAOUT8 ;
wire \mac_mult8~DATAOUT9 ;
wire \mac_mult8~DATAOUT10 ;
wire \mac_mult8~DATAOUT11 ;
wire \mac_mult8~DATAOUT12 ;
wire \mac_mult8~DATAOUT13 ;
wire \mac_mult8~DATAOUT14 ;
wire \mac_mult8~DATAOUT15 ;

wire [35:0] mac_out9_DATAOUT_bus;
wire [35:0] mac_mult8_DATAOUT_bus;

assign mac_out91 = mac_out9_DATAOUT_bus[0];
assign mac_out92 = mac_out9_DATAOUT_bus[1];
assign mac_out93 = mac_out9_DATAOUT_bus[2];
assign mac_out94 = mac_out9_DATAOUT_bus[3];
assign mac_out95 = mac_out9_DATAOUT_bus[4];
assign mac_out96 = mac_out9_DATAOUT_bus[5];
assign mac_out97 = mac_out9_DATAOUT_bus[6];
assign mac_out98 = mac_out9_DATAOUT_bus[7];
assign mac_out99 = mac_out9_DATAOUT_bus[8];
assign mac_out910 = mac_out9_DATAOUT_bus[9];
assign mac_out911 = mac_out9_DATAOUT_bus[10];
assign mac_out912 = mac_out9_DATAOUT_bus[11];
assign mac_out913 = mac_out9_DATAOUT_bus[12];
assign mac_out914 = mac_out9_DATAOUT_bus[13];
assign mac_out915 = mac_out9_DATAOUT_bus[14];
assign mac_out916 = mac_out9_DATAOUT_bus[15];

assign \mac_mult8~dataout  = mac_mult8_DATAOUT_bus[0];
assign \mac_mult8~DATAOUT1  = mac_mult8_DATAOUT_bus[1];
assign \mac_mult8~DATAOUT2  = mac_mult8_DATAOUT_bus[2];
assign \mac_mult8~DATAOUT3  = mac_mult8_DATAOUT_bus[3];
assign \mac_mult8~DATAOUT4  = mac_mult8_DATAOUT_bus[4];
assign \mac_mult8~DATAOUT5  = mac_mult8_DATAOUT_bus[5];
assign \mac_mult8~DATAOUT6  = mac_mult8_DATAOUT_bus[6];
assign \mac_mult8~DATAOUT7  = mac_mult8_DATAOUT_bus[7];
assign \mac_mult8~DATAOUT8  = mac_mult8_DATAOUT_bus[8];
assign \mac_mult8~DATAOUT9  = mac_mult8_DATAOUT_bus[9];
assign \mac_mult8~DATAOUT10  = mac_mult8_DATAOUT_bus[10];
assign \mac_mult8~DATAOUT11  = mac_mult8_DATAOUT_bus[11];
assign \mac_mult8~DATAOUT12  = mac_mult8_DATAOUT_bus[12];
assign \mac_mult8~DATAOUT13  = mac_mult8_DATAOUT_bus[13];
assign \mac_mult8~DATAOUT14  = mac_mult8_DATAOUT_bus[14];
assign \mac_mult8~DATAOUT15  = mac_mult8_DATAOUT_bus[15];

cycloneiv_mac_out mac_out9(
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\mac_mult8~DATAOUT15 ,\mac_mult8~DATAOUT14 ,\mac_mult8~DATAOUT13 ,\mac_mult8~DATAOUT12 ,\mac_mult8~DATAOUT11 ,\mac_mult8~DATAOUT10 ,\mac_mult8~DATAOUT9 ,\mac_mult8~DATAOUT8 ,\mac_mult8~DATAOUT7 ,
\mac_mult8~DATAOUT6 ,\mac_mult8~DATAOUT5 ,\mac_mult8~DATAOUT4 ,\mac_mult8~DATAOUT3 ,\mac_mult8~DATAOUT2 ,\mac_mult8~DATAOUT1 ,\mac_mult8~dataout }),
	.dataout(mac_out9_DATAOUT_bus));
defparam mac_out9.dataa_width = 16;
defparam mac_out9.output_clock = "0";

cycloneiv_mac_mult mac_mult8(
	.signa(vcc),
	.signb(vcc),
	.clk(clock[0]),
	.aclr(!aclr[0]),
	.ena(ena[0]),
	.dataa({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,dataa[7],dataa[6],dataa[5],dataa[4],dataa[3],dataa[2],dataa[1],dataa[0]}),
	.datab({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,datab[7],datab[6],datab[5],datab[4],datab[3],datab[2],datab[1],datab[0]}),
	.dataout(mac_mult8_DATAOUT_bus));
defparam mac_mult8.dataa_clock = "0";
defparam mac_mult8.dataa_width = 8;
defparam mac_mult8.datab_clock = "0";
defparam mac_mult8.datab_width = 8;
defparam mac_mult8.signa_clock = "none";
defparam mac_mult8.signb_clock = "none";

endmodule

module ifft_8p_auk_dspip_r22sdf_counter_3 (
	stg_valid_next,
	curr_pwr_2_s,
	out_enable,
	stg_sop_next,
	control_s_1,
	control_s_2,
	control_s_0,
	stg_control_next_1,
	stg_control_next_2,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
input 	stg_valid_next;
input 	curr_pwr_2_s;
input 	out_enable;
input 	stg_sop_next;
output 	control_s_1;
output 	control_s_2;
output 	control_s_0;
input 	stg_control_next_1;
input 	stg_control_next_2;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \control_s~0_combout ;
wire \counter_p~0_combout ;
wire \control_s~1_combout ;
wire \control_s~2_combout ;
wire \control_s~3_combout ;


dffeas \control_s[1] (
	.clk(clk),
	.d(\control_s~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_p~0_combout ),
	.q(control_s_1),
	.prn(vcc));
defparam \control_s[1] .is_wysiwyg = "true";
defparam \control_s[1] .power_up = "low";

dffeas \control_s[2] (
	.clk(clk),
	.d(\control_s~2_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_p~0_combout ),
	.q(control_s_2),
	.prn(vcc));
defparam \control_s[2] .is_wysiwyg = "true";
defparam \control_s[2] .power_up = "low";

dffeas \control_s[0] (
	.clk(clk),
	.d(\control_s~3_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\counter_p~0_combout ),
	.q(control_s_0),
	.prn(vcc));
defparam \control_s[0] .is_wysiwyg = "true";
defparam \control_s[0] .power_up = "low";

cycloneiv_lcell_comb \control_s~0 (
	.dataa(control_s_1),
	.datab(control_s_0),
	.datac(stg_sop_next),
	.datad(stg_control_next_1),
	.cin(gnd),
	.combout(\control_s~0_combout ),
	.cout());
defparam \control_s~0 .lut_mask = 16'h96FF;
defparam \control_s~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \counter_p~0 (
	.dataa(curr_pwr_2_s),
	.datab(stg_valid_next),
	.datac(gnd),
	.datad(out_enable),
	.cin(gnd),
	.combout(\counter_p~0_combout ),
	.cout());
defparam \counter_p~0 .lut_mask = 16'hFFEE;
defparam \counter_p~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~1 (
	.dataa(control_s_2),
	.datab(control_s_1),
	.datac(control_s_0),
	.datad(stg_sop_next),
	.cin(gnd),
	.combout(\control_s~1_combout ),
	.cout());
defparam \control_s~1 .lut_mask = 16'h96FF;
defparam \control_s~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~2 (
	.dataa(\control_s~1_combout ),
	.datab(stg_sop_next),
	.datac(stg_control_next_1),
	.datad(stg_control_next_2),
	.cin(gnd),
	.combout(\control_s~2_combout ),
	.cout());
defparam \control_s~2 .lut_mask = 16'hEFFE;
defparam \control_s~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \control_s~3 (
	.dataa(stg_sop_next),
	.datab(control_s_0),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\control_s~3_combout ),
	.cout());
defparam \control_s~3 .lut_mask = 16'h7777;
defparam \control_s~3 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_roundsat (
	dataout_2,
	dataout_1,
	dataout_0,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	out_stall_d,
	sop,
	out_valid_s,
	out_sop_d_2,
	conv_round_3OR_accu,
	NONA10_C_Mult_Archsgen_small_multimag_result9,
	NONA10_C_Mult_Archsgen_small_multimag_result8,
	NONA10_C_Mult_Archsgen_small_multimag_result7,
	NONA10_C_Mult_Archsgen_small_multimag_result6,
	NONA10_C_Mult_Archsgen_small_multimag_result3,
	NONA10_C_Mult_Archsgen_small_multimag_result4,
	NONA10_C_Mult_Archsgen_small_multimag_result5,
	NONA10_C_Mult_Archsgen_small_multimag_result0,
	NONA10_C_Mult_Archsgen_small_multimag_result1,
	NONA10_C_Mult_Archsgen_small_multimag_result2,
	NONA10_C_Mult_Archsgen_small_multimag_result10,
	NONA10_C_Mult_Archsgen_small_multimag_result11,
	NONA10_C_Mult_Archsgen_small_multimag_result12,
	NONA10_C_Mult_Archsgen_small_multimag_result13,
	NONA10_C_Mult_Archsgen_small_multimag_result14,
	NONA10_C_Mult_Archsgen_small_multimag_result15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dataout_2;
output 	dataout_1;
output 	dataout_0;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
input 	out_stall_d;
input 	sop;
input 	out_valid_s;
input 	out_sop_d_2;
output 	conv_round_3OR_accu;
input 	NONA10_C_Mult_Archsgen_small_multimag_result9;
input 	NONA10_C_Mult_Archsgen_small_multimag_result8;
input 	NONA10_C_Mult_Archsgen_small_multimag_result7;
input 	NONA10_C_Mult_Archsgen_small_multimag_result6;
input 	NONA10_C_Mult_Archsgen_small_multimag_result3;
input 	NONA10_C_Mult_Archsgen_small_multimag_result4;
input 	NONA10_C_Mult_Archsgen_small_multimag_result5;
input 	NONA10_C_Mult_Archsgen_small_multimag_result0;
input 	NONA10_C_Mult_Archsgen_small_multimag_result1;
input 	NONA10_C_Mult_Archsgen_small_multimag_result2;
input 	NONA10_C_Mult_Archsgen_small_multimag_result10;
input 	NONA10_C_Mult_Archsgen_small_multimag_result11;
input 	NONA10_C_Mult_Archsgen_small_multimag_result12;
input 	NONA10_C_Mult_Archsgen_small_multimag_result13;
input 	NONA10_C_Mult_Archsgen_small_multimag_result14;
input 	NONA10_C_Mult_Archsgen_small_multimag_result15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \datareg~0_combout ;
wire \conv_round_3:datareg[9]~q ;
wire \conv_round_3:datareg_2[9]~q ;
wire \datareg~1_combout ;
wire \conv_round_3:datareg[8]~q ;
wire \conv_round_3:datareg_2[8]~q ;
wire \LSB~0_combout ;
wire \conv_round_3:LSB~q ;
wire \conv_round_3:datareg_2[7]~q ;
wire \RB~0_combout ;
wire \conv_round_3:RB~q ;
wire \RB_R~0_combout ;
wire \conv_round_3:RB_R~q ;
wire \OR_Temp_2~0_combout ;
wire \conv_round_3:OR_accu_2~q ;
wire \OR_Temp_1~0_combout ;
wire \conv_round_3:OR_accu_1~q ;
wire \OR_accu~0_combout ;
wire \conv_round_3:OR_accu~q ;
wire \LSB_R~0_combout ;
wire \conv_round_3:LSB_R~q ;
wire \conv_round_p2~0_combout ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~2_combout ;
wire \Add0~0_combout ;
wire \datareg~2_combout ;
wire \conv_round_3:datareg[10]~q ;
wire \conv_round_3:datareg_2[10]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \datareg~3_combout ;
wire \conv_round_3:datareg[11]~q ;
wire \conv_round_3:datareg_2[11]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \datareg~4_combout ;
wire \conv_round_3:datareg[12]~q ;
wire \conv_round_3:datareg_2[12]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \datareg~5_combout ;
wire \conv_round_3:datareg[13]~q ;
wire \conv_round_3:datareg_2[13]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \datareg~6_combout ;
wire \conv_round_3:datareg[14]~q ;
wire \conv_round_3:datareg_2[14]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \datareg~7_combout ;
wire \conv_round_3:datareg[15]~q ;
wire \conv_round_3:datareg_2[15]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;


dffeas \dataout[2] (
	.clk(clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_2),
	.prn(vcc));
defparam \dataout[2] .is_wysiwyg = "true";
defparam \dataout[2] .power_up = "low";

dffeas \dataout[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_1),
	.prn(vcc));
defparam \dataout[1] .is_wysiwyg = "true";
defparam \dataout[1] .power_up = "low";

dffeas \dataout[0] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_0),
	.prn(vcc));
defparam \dataout[0] .is_wysiwyg = "true";
defparam \dataout[0] .power_up = "low";

dffeas \dataout[3] (
	.clk(clk),
	.d(\Add0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_3),
	.prn(vcc));
defparam \dataout[3] .is_wysiwyg = "true";
defparam \dataout[3] .power_up = "low";

dffeas \dataout[4] (
	.clk(clk),
	.d(\Add0~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_4),
	.prn(vcc));
defparam \dataout[4] .is_wysiwyg = "true";
defparam \dataout[4] .power_up = "low";

dffeas \dataout[5] (
	.clk(clk),
	.d(\Add0~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_5),
	.prn(vcc));
defparam \dataout[5] .is_wysiwyg = "true";
defparam \dataout[5] .power_up = "low";

dffeas \dataout[6] (
	.clk(clk),
	.d(\Add0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_6),
	.prn(vcc));
defparam \dataout[6] .is_wysiwyg = "true";
defparam \dataout[6] .power_up = "low";

dffeas \dataout[7] (
	.clk(clk),
	.d(\Add0~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_7),
	.prn(vcc));
defparam \dataout[7] .is_wysiwyg = "true";
defparam \dataout[7] .power_up = "low";

dffeas \dataout[8] (
	.clk(clk),
	.d(\Add0~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_8),
	.prn(vcc));
defparam \dataout[8] .is_wysiwyg = "true";
defparam \dataout[8] .power_up = "low";

cycloneiv_lcell_comb \conv_round_3:OR_accu~0 (
	.dataa(reset_n),
	.datab(out_valid_s),
	.datac(sop),
	.datad(out_stall_d),
	.cin(gnd),
	.combout(conv_round_3OR_accu),
	.cout());
defparam \conv_round_3:OR_accu~0 .lut_mask = 16'hACFF;
defparam \conv_round_3:OR_accu~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \datareg~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~0_combout ),
	.cout());
defparam \datareg~0 .lut_mask = 16'hEEEE;
defparam \datareg~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[9] (
	.clk(clk),
	.d(\datareg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[9]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[9] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[9] .power_up = "low";

dffeas \conv_round_3:datareg_2[9] (
	.clk(clk),
	.d(\conv_round_3:datareg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[9]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[9] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[9] .power_up = "low";

cycloneiv_lcell_comb \datareg~1 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~1_combout ),
	.cout());
defparam \datareg~1 .lut_mask = 16'hEEEE;
defparam \datareg~1 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[8] (
	.clk(clk),
	.d(\datareg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[8]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[8] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[8] .power_up = "low";

dffeas \conv_round_3:datareg_2[8] (
	.clk(clk),
	.d(\conv_round_3:datareg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[8]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[8] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[8] .power_up = "low";

cycloneiv_lcell_comb \LSB~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LSB~0_combout ),
	.cout());
defparam \LSB~0 .lut_mask = 16'hEEEE;
defparam \LSB~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:LSB (
	.clk(clk),
	.d(\LSB~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:LSB~q ),
	.prn(vcc));
defparam \conv_round_3:LSB .is_wysiwyg = "true";
defparam \conv_round_3:LSB .power_up = "low";

dffeas \conv_round_3:datareg_2[7] (
	.clk(clk),
	.d(\conv_round_3:LSB~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[7]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[7] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[7] .power_up = "low";

cycloneiv_lcell_comb \RB~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\RB~0_combout ),
	.cout());
defparam \RB~0 .lut_mask = 16'hEEEE;
defparam \RB~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:RB (
	.clk(clk),
	.d(\RB~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:RB~q ),
	.prn(vcc));
defparam \conv_round_3:RB .is_wysiwyg = "true";
defparam \conv_round_3:RB .power_up = "low";

cycloneiv_lcell_comb \RB_R~0 (
	.dataa(reset_n),
	.datab(\conv_round_3:RB~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\RB_R~0_combout ),
	.cout());
defparam \RB_R~0 .lut_mask = 16'hEEEE;
defparam \RB_R~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:RB_R (
	.clk(clk),
	.d(\RB_R~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:RB_R~q ),
	.prn(vcc));
defparam \conv_round_3:RB_R .is_wysiwyg = "true";
defparam \conv_round_3:RB_R .power_up = "low";

cycloneiv_lcell_comb \OR_Temp_2~0 (
	.dataa(NONA10_C_Mult_Archsgen_small_multimag_result3),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result4),
	.datac(NONA10_C_Mult_Archsgen_small_multimag_result5),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_Temp_2~0_combout ),
	.cout());
defparam \OR_Temp_2~0 .lut_mask = 16'hFEFE;
defparam \OR_Temp_2~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu_2 (
	.clk(clk),
	.d(\OR_Temp_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:OR_accu_2~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu_2 .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu_2 .power_up = "low";

cycloneiv_lcell_comb \OR_Temp_1~0 (
	.dataa(NONA10_C_Mult_Archsgen_small_multimag_result0),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result1),
	.datac(NONA10_C_Mult_Archsgen_small_multimag_result2),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_Temp_1~0_combout ),
	.cout());
defparam \OR_Temp_1~0 .lut_mask = 16'hFEFE;
defparam \OR_Temp_1~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu_1 (
	.clk(clk),
	.d(\OR_Temp_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:OR_accu_1~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu_1 .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu_1 .power_up = "low";

cycloneiv_lcell_comb \OR_accu~0 (
	.dataa(\conv_round_3:OR_accu_2~q ),
	.datab(\conv_round_3:OR_accu_1~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_accu~0_combout ),
	.cout());
defparam \OR_accu~0 .lut_mask = 16'hEEEE;
defparam \OR_accu~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu (
	.clk(clk),
	.d(\OR_accu~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:OR_accu~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu .power_up = "low";

cycloneiv_lcell_comb \LSB_R~0 (
	.dataa(reset_n),
	.datab(\conv_round_3:LSB~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LSB_R~0_combout ),
	.cout());
defparam \LSB_R~0 .lut_mask = 16'hEEEE;
defparam \LSB_R~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:LSB_R (
	.clk(clk),
	.d(\LSB_R~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:LSB_R~q ),
	.prn(vcc));
defparam \conv_round_3:LSB_R .is_wysiwyg = "true";
defparam \conv_round_3:LSB_R .power_up = "low";

cycloneiv_lcell_comb \conv_round_p2~0 (
	.dataa(\conv_round_3:RB_R~q ),
	.datab(\conv_round_3:OR_accu~q ),
	.datac(\conv_round_3:LSB_R~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\conv_round_p2~0_combout ),
	.cout());
defparam \conv_round_p2~0 .lut_mask = 16'hFEFE;
defparam \conv_round_p2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~0 (
	.dataa(\conv_round_3:datareg_2[7]~q ),
	.datab(\conv_round_p2~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h66EE;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~2 (
	.dataa(\conv_round_3:datareg_2[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add0~4 (
	.dataa(\conv_round_3:datareg_2[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~2 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~2_combout ),
	.cout());
defparam \datareg~2 .lut_mask = 16'hEEEE;
defparam \datareg~2 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[10] (
	.clk(clk),
	.d(\datareg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[10]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[10] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[10] .power_up = "low";

dffeas \conv_round_3:datareg_2[10] (
	.clk(clk),
	.d(\conv_round_3:datareg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[10]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[10] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[10] .power_up = "low";

cycloneiv_lcell_comb \Add0~6 (
	.dataa(\conv_round_3:datareg_2[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~3 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~3_combout ),
	.cout());
defparam \datareg~3 .lut_mask = 16'hEEEE;
defparam \datareg~3 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[11] (
	.clk(clk),
	.d(\datareg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[11]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[11] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[11] .power_up = "low";

dffeas \conv_round_3:datareg_2[11] (
	.clk(clk),
	.d(\conv_round_3:datareg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[11]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[11] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[11] .power_up = "low";

cycloneiv_lcell_comb \Add0~8 (
	.dataa(\conv_round_3:datareg_2[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~4 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~4_combout ),
	.cout());
defparam \datareg~4 .lut_mask = 16'hEEEE;
defparam \datareg~4 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[12] (
	.clk(clk),
	.d(\datareg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[12]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[12] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[12] .power_up = "low";

dffeas \conv_round_3:datareg_2[12] (
	.clk(clk),
	.d(\conv_round_3:datareg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[12]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[12] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[12] .power_up = "low";

cycloneiv_lcell_comb \Add0~10 (
	.dataa(\conv_round_3:datareg_2[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~5 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~5_combout ),
	.cout());
defparam \datareg~5 .lut_mask = 16'hEEEE;
defparam \datareg~5 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[13] (
	.clk(clk),
	.d(\datareg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[13]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[13] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[13] .power_up = "low";

dffeas \conv_round_3:datareg_2[13] (
	.clk(clk),
	.d(\conv_round_3:datareg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[13]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[13] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[13] .power_up = "low";

cycloneiv_lcell_comb \Add0~12 (
	.dataa(\conv_round_3:datareg_2[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~6 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~6_combout ),
	.cout());
defparam \datareg~6 .lut_mask = 16'hEEEE;
defparam \datareg~6 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[14] (
	.clk(clk),
	.d(\datareg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[14]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[14] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[14] .power_up = "low";

dffeas \conv_round_3:datareg_2[14] (
	.clk(clk),
	.d(\conv_round_3:datareg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[14]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[14] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[14] .power_up = "low";

cycloneiv_lcell_comb \Add0~14 (
	.dataa(\conv_round_3:datareg_2[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~7 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multimag_result15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~7_combout ),
	.cout());
defparam \datareg~7 .lut_mask = 16'hEEEE;
defparam \datareg~7 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[15] (
	.clk(clk),
	.d(\datareg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[15]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[15] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[15] .power_up = "low";

dffeas \conv_round_3:datareg_2[15] (
	.clk(clk),
	.d(\conv_round_3:datareg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(conv_round_3OR_accu),
	.q(\conv_round_3:datareg_2[15]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[15] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[15] .power_up = "low";

cycloneiv_lcell_comb \Add0~16 (
	.dataa(\conv_round_3:datareg_2[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout());
defparam \Add0~16 .lut_mask = 16'h5A5A;
defparam \Add0~16 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_roundsat_1 (
	dataout_2,
	dataout_1,
	dataout_0,
	dataout_3,
	dataout_4,
	dataout_5,
	dataout_6,
	dataout_7,
	dataout_8,
	out_sop_d_2,
	reset,
	NONA10_C_Mult_Archsgen_small_multreal_result9,
	NONA10_C_Mult_Archsgen_small_multreal_result8,
	NONA10_C_Mult_Archsgen_small_multreal_result7,
	NONA10_C_Mult_Archsgen_small_multreal_result6,
	NONA10_C_Mult_Archsgen_small_multreal_result3,
	NONA10_C_Mult_Archsgen_small_multreal_result4,
	NONA10_C_Mult_Archsgen_small_multreal_result5,
	NONA10_C_Mult_Archsgen_small_multreal_result0,
	NONA10_C_Mult_Archsgen_small_multreal_result1,
	NONA10_C_Mult_Archsgen_small_multreal_result2,
	NONA10_C_Mult_Archsgen_small_multreal_result10,
	NONA10_C_Mult_Archsgen_small_multreal_result11,
	NONA10_C_Mult_Archsgen_small_multreal_result12,
	NONA10_C_Mult_Archsgen_small_multreal_result13,
	NONA10_C_Mult_Archsgen_small_multreal_result14,
	NONA10_C_Mult_Archsgen_small_multreal_result15,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	dataout_2;
output 	dataout_1;
output 	dataout_0;
output 	dataout_3;
output 	dataout_4;
output 	dataout_5;
output 	dataout_6;
output 	dataout_7;
output 	dataout_8;
input 	out_sop_d_2;
input 	reset;
input 	NONA10_C_Mult_Archsgen_small_multreal_result9;
input 	NONA10_C_Mult_Archsgen_small_multreal_result8;
input 	NONA10_C_Mult_Archsgen_small_multreal_result7;
input 	NONA10_C_Mult_Archsgen_small_multreal_result6;
input 	NONA10_C_Mult_Archsgen_small_multreal_result3;
input 	NONA10_C_Mult_Archsgen_small_multreal_result4;
input 	NONA10_C_Mult_Archsgen_small_multreal_result5;
input 	NONA10_C_Mult_Archsgen_small_multreal_result0;
input 	NONA10_C_Mult_Archsgen_small_multreal_result1;
input 	NONA10_C_Mult_Archsgen_small_multreal_result2;
input 	NONA10_C_Mult_Archsgen_small_multreal_result10;
input 	NONA10_C_Mult_Archsgen_small_multreal_result11;
input 	NONA10_C_Mult_Archsgen_small_multreal_result12;
input 	NONA10_C_Mult_Archsgen_small_multreal_result13;
input 	NONA10_C_Mult_Archsgen_small_multreal_result14;
input 	NONA10_C_Mult_Archsgen_small_multreal_result15;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \datareg~0_combout ;
wire \conv_round_3:datareg[9]~q ;
wire \conv_round_3:datareg_2[9]~q ;
wire \datareg~1_combout ;
wire \conv_round_3:datareg[8]~q ;
wire \conv_round_3:datareg_2[8]~q ;
wire \LSB~0_combout ;
wire \conv_round_3:LSB~q ;
wire \conv_round_3:datareg_2[7]~q ;
wire \RB~0_combout ;
wire \conv_round_3:RB~q ;
wire \RB_R~0_combout ;
wire \conv_round_3:RB_R~q ;
wire \OR_Temp_2~0_combout ;
wire \conv_round_3:OR_accu_2~q ;
wire \OR_Temp_1~0_combout ;
wire \conv_round_3:OR_accu_1~q ;
wire \OR_accu~0_combout ;
wire \conv_round_3:OR_accu~q ;
wire \LSB_R~0_combout ;
wire \conv_round_3:LSB_R~q ;
wire \conv_round_p2~0_combout ;
wire \Add0~1 ;
wire \Add0~3 ;
wire \Add0~4_combout ;
wire \Add0~2_combout ;
wire \Add0~0_combout ;
wire \datareg~2_combout ;
wire \conv_round_3:datareg[10]~q ;
wire \conv_round_3:datareg_2[10]~q ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \datareg~3_combout ;
wire \conv_round_3:datareg[11]~q ;
wire \conv_round_3:datareg_2[11]~q ;
wire \Add0~7 ;
wire \Add0~8_combout ;
wire \datareg~4_combout ;
wire \conv_round_3:datareg[12]~q ;
wire \conv_round_3:datareg_2[12]~q ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \datareg~5_combout ;
wire \conv_round_3:datareg[13]~q ;
wire \conv_round_3:datareg_2[13]~q ;
wire \Add0~11 ;
wire \Add0~12_combout ;
wire \datareg~6_combout ;
wire \conv_round_3:datareg[14]~q ;
wire \conv_round_3:datareg_2[14]~q ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \datareg~7_combout ;
wire \conv_round_3:datareg[15]~q ;
wire \conv_round_3:datareg_2[15]~q ;
wire \Add0~15 ;
wire \Add0~16_combout ;


dffeas \dataout[2] (
	.clk(clk),
	.d(\Add0~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_2),
	.prn(vcc));
defparam \dataout[2] .is_wysiwyg = "true";
defparam \dataout[2] .power_up = "low";

dffeas \dataout[1] (
	.clk(clk),
	.d(\Add0~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_1),
	.prn(vcc));
defparam \dataout[1] .is_wysiwyg = "true";
defparam \dataout[1] .power_up = "low";

dffeas \dataout[0] (
	.clk(clk),
	.d(\Add0~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_0),
	.prn(vcc));
defparam \dataout[0] .is_wysiwyg = "true";
defparam \dataout[0] .power_up = "low";

dffeas \dataout[3] (
	.clk(clk),
	.d(\Add0~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_3),
	.prn(vcc));
defparam \dataout[3] .is_wysiwyg = "true";
defparam \dataout[3] .power_up = "low";

dffeas \dataout[4] (
	.clk(clk),
	.d(\Add0~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_4),
	.prn(vcc));
defparam \dataout[4] .is_wysiwyg = "true";
defparam \dataout[4] .power_up = "low";

dffeas \dataout[5] (
	.clk(clk),
	.d(\Add0~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_5),
	.prn(vcc));
defparam \dataout[5] .is_wysiwyg = "true";
defparam \dataout[5] .power_up = "low";

dffeas \dataout[6] (
	.clk(clk),
	.d(\Add0~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_6),
	.prn(vcc));
defparam \dataout[6] .is_wysiwyg = "true";
defparam \dataout[6] .power_up = "low";

dffeas \dataout[7] (
	.clk(clk),
	.d(\Add0~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_7),
	.prn(vcc));
defparam \dataout[7] .is_wysiwyg = "true";
defparam \dataout[7] .power_up = "low";

dffeas \dataout[8] (
	.clk(clk),
	.d(\Add0~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(dataout_8),
	.prn(vcc));
defparam \dataout[8] .is_wysiwyg = "true";
defparam \dataout[8] .power_up = "low";

cycloneiv_lcell_comb \datareg~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result9),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~0_combout ),
	.cout());
defparam \datareg~0 .lut_mask = 16'hEEEE;
defparam \datareg~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[9] (
	.clk(clk),
	.d(\datareg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[9]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[9] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[9] .power_up = "low";

dffeas \conv_round_3:datareg_2[9] (
	.clk(clk),
	.d(\conv_round_3:datareg[9]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[9]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[9] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[9] .power_up = "low";

cycloneiv_lcell_comb \datareg~1 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result8),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~1_combout ),
	.cout());
defparam \datareg~1 .lut_mask = 16'hEEEE;
defparam \datareg~1 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[8] (
	.clk(clk),
	.d(\datareg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[8]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[8] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[8] .power_up = "low";

dffeas \conv_round_3:datareg_2[8] (
	.clk(clk),
	.d(\conv_round_3:datareg[8]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[8]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[8] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[8] .power_up = "low";

cycloneiv_lcell_comb \LSB~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result7),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LSB~0_combout ),
	.cout());
defparam \LSB~0 .lut_mask = 16'hEEEE;
defparam \LSB~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:LSB (
	.clk(clk),
	.d(\LSB~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:LSB~q ),
	.prn(vcc));
defparam \conv_round_3:LSB .is_wysiwyg = "true";
defparam \conv_round_3:LSB .power_up = "low";

dffeas \conv_round_3:datareg_2[7] (
	.clk(clk),
	.d(\conv_round_3:LSB~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[7]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[7] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[7] .power_up = "low";

cycloneiv_lcell_comb \RB~0 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result6),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\RB~0_combout ),
	.cout());
defparam \RB~0 .lut_mask = 16'hEEEE;
defparam \RB~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:RB (
	.clk(clk),
	.d(\RB~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:RB~q ),
	.prn(vcc));
defparam \conv_round_3:RB .is_wysiwyg = "true";
defparam \conv_round_3:RB .power_up = "low";

cycloneiv_lcell_comb \RB_R~0 (
	.dataa(reset_n),
	.datab(\conv_round_3:RB~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\RB_R~0_combout ),
	.cout());
defparam \RB_R~0 .lut_mask = 16'hEEEE;
defparam \RB_R~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:RB_R (
	.clk(clk),
	.d(\RB_R~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:RB_R~q ),
	.prn(vcc));
defparam \conv_round_3:RB_R .is_wysiwyg = "true";
defparam \conv_round_3:RB_R .power_up = "low";

cycloneiv_lcell_comb \OR_Temp_2~0 (
	.dataa(NONA10_C_Mult_Archsgen_small_multreal_result3),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result4),
	.datac(NONA10_C_Mult_Archsgen_small_multreal_result5),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_Temp_2~0_combout ),
	.cout());
defparam \OR_Temp_2~0 .lut_mask = 16'hFEFE;
defparam \OR_Temp_2~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu_2 (
	.clk(clk),
	.d(\OR_Temp_2~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:OR_accu_2~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu_2 .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu_2 .power_up = "low";

cycloneiv_lcell_comb \OR_Temp_1~0 (
	.dataa(NONA10_C_Mult_Archsgen_small_multreal_result0),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result1),
	.datac(NONA10_C_Mult_Archsgen_small_multreal_result2),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_Temp_1~0_combout ),
	.cout());
defparam \OR_Temp_1~0 .lut_mask = 16'hFEFE;
defparam \OR_Temp_1~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu_1 (
	.clk(clk),
	.d(\OR_Temp_1~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!reset_n),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:OR_accu_1~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu_1 .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu_1 .power_up = "low";

cycloneiv_lcell_comb \OR_accu~0 (
	.dataa(\conv_round_3:OR_accu_2~q ),
	.datab(\conv_round_3:OR_accu_1~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\OR_accu~0_combout ),
	.cout());
defparam \OR_accu~0 .lut_mask = 16'hEEEE;
defparam \OR_accu~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:OR_accu (
	.clk(clk),
	.d(\OR_accu~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:OR_accu~q ),
	.prn(vcc));
defparam \conv_round_3:OR_accu .is_wysiwyg = "true";
defparam \conv_round_3:OR_accu .power_up = "low";

cycloneiv_lcell_comb \LSB_R~0 (
	.dataa(reset_n),
	.datab(\conv_round_3:LSB~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\LSB_R~0_combout ),
	.cout());
defparam \LSB_R~0 .lut_mask = 16'hEEEE;
defparam \LSB_R~0 .sum_lutc_input = "datac";

dffeas \conv_round_3:LSB_R (
	.clk(clk),
	.d(\LSB_R~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:LSB_R~q ),
	.prn(vcc));
defparam \conv_round_3:LSB_R .is_wysiwyg = "true";
defparam \conv_round_3:LSB_R .power_up = "low";

cycloneiv_lcell_comb \conv_round_p2~0 (
	.dataa(\conv_round_3:RB_R~q ),
	.datab(\conv_round_3:OR_accu~q ),
	.datac(\conv_round_3:LSB_R~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\conv_round_p2~0_combout ),
	.cout());
defparam \conv_round_p2~0 .lut_mask = 16'hFEFE;
defparam \conv_round_p2~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~0 (
	.dataa(\conv_round_3:datareg_2[7]~q ),
	.datab(\conv_round_p2~0_combout ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
defparam \Add0~0 .lut_mask = 16'h66EE;
defparam \Add0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add0~2 (
	.dataa(\conv_round_3:datareg_2[8]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
defparam \Add0~2 .lut_mask = 16'h5A5F;
defparam \Add0~2 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add0~4 (
	.dataa(\conv_round_3:datareg_2[9]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
defparam \Add0~4 .lut_mask = 16'h5AAF;
defparam \Add0~4 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~2 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result10),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~2_combout ),
	.cout());
defparam \datareg~2 .lut_mask = 16'hEEEE;
defparam \datareg~2 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[10] (
	.clk(clk),
	.d(\datareg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[10]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[10] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[10] .power_up = "low";

dffeas \conv_round_3:datareg_2[10] (
	.clk(clk),
	.d(\conv_round_3:datareg[10]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[10]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[10] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[10] .power_up = "low";

cycloneiv_lcell_comb \Add0~6 (
	.dataa(\conv_round_3:datareg_2[10]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
defparam \Add0~6 .lut_mask = 16'h5A5F;
defparam \Add0~6 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~3 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result11),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~3_combout ),
	.cout());
defparam \datareg~3 .lut_mask = 16'hEEEE;
defparam \datareg~3 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[11] (
	.clk(clk),
	.d(\datareg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[11]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[11] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[11] .power_up = "low";

dffeas \conv_round_3:datareg_2[11] (
	.clk(clk),
	.d(\conv_round_3:datareg[11]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[11]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[11] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[11] .power_up = "low";

cycloneiv_lcell_comb \Add0~8 (
	.dataa(\conv_round_3:datareg_2[11]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
defparam \Add0~8 .lut_mask = 16'h5AAF;
defparam \Add0~8 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~4 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result12),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~4_combout ),
	.cout());
defparam \datareg~4 .lut_mask = 16'hEEEE;
defparam \datareg~4 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[12] (
	.clk(clk),
	.d(\datareg~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[12]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[12] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[12] .power_up = "low";

dffeas \conv_round_3:datareg_2[12] (
	.clk(clk),
	.d(\conv_round_3:datareg[12]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[12]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[12] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[12] .power_up = "low";

cycloneiv_lcell_comb \Add0~10 (
	.dataa(\conv_round_3:datareg_2[12]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
defparam \Add0~10 .lut_mask = 16'h5A5F;
defparam \Add0~10 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~5 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result13),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~5_combout ),
	.cout());
defparam \datareg~5 .lut_mask = 16'hEEEE;
defparam \datareg~5 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[13] (
	.clk(clk),
	.d(\datareg~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[13]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[13] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[13] .power_up = "low";

dffeas \conv_round_3:datareg_2[13] (
	.clk(clk),
	.d(\conv_round_3:datareg[13]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[13]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[13] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[13] .power_up = "low";

cycloneiv_lcell_comb \Add0~12 (
	.dataa(\conv_round_3:datareg_2[13]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
defparam \Add0~12 .lut_mask = 16'h5AAF;
defparam \Add0~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~6 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result14),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~6_combout ),
	.cout());
defparam \datareg~6 .lut_mask = 16'hEEEE;
defparam \datareg~6 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[14] (
	.clk(clk),
	.d(\datareg~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[14]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[14] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[14] .power_up = "low";

dffeas \conv_round_3:datareg_2[14] (
	.clk(clk),
	.d(\conv_round_3:datareg[14]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[14]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[14] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[14] .power_up = "low";

cycloneiv_lcell_comb \Add0~14 (
	.dataa(\conv_round_3:datareg_2[14]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
defparam \Add0~14 .lut_mask = 16'h5A5F;
defparam \Add0~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \datareg~7 (
	.dataa(reset_n),
	.datab(NONA10_C_Mult_Archsgen_small_multreal_result15),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\datareg~7_combout ),
	.cout());
defparam \datareg~7 .lut_mask = 16'hEEEE;
defparam \datareg~7 .sum_lutc_input = "datac";

dffeas \conv_round_3:datareg[15] (
	.clk(clk),
	.d(\datareg~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_sop_d_2),
	.q(\conv_round_3:datareg[15]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg[15] .is_wysiwyg = "true";
defparam \conv_round_3:datareg[15] .power_up = "low";

dffeas \conv_round_3:datareg_2[15] (
	.clk(clk),
	.d(\conv_round_3:datareg[15]~q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(reset),
	.q(\conv_round_3:datareg_2[15]~q ),
	.prn(vcc));
defparam \conv_round_3:datareg_2[15] .is_wysiwyg = "true";
defparam \conv_round_3:datareg_2[15] .power_up = "low";

cycloneiv_lcell_comb \Add0~16 (
	.dataa(\conv_round_3:datareg_2[15]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout());
defparam \Add0~16 .lut_mask = 16'h5A5A;
defparam \Add0~16 .sum_lutc_input = "cin";

endmodule

module ifft_8p_auk_dspip_r22sdf_stg_pipe (
	stg_imag_next_0,
	stg_real_next_0,
	stg_imag_next_1,
	stg_real_next_1,
	stg_imag_next_2,
	stg_real_next_2,
	stg_imag_next_3,
	stg_real_next_3,
	stg_imag_next_4,
	stg_real_next_4,
	stg_imag_next_5,
	stg_real_next_5,
	stg_imag_next_6,
	stg_real_next_6,
	stg_imag_next_7,
	stg_real_next_7,
	stg_imag_next_01,
	out_imag_2,
	stg_real_next_01,
	out_real_2,
	stg_imag_next_11,
	out_imag_3,
	stg_real_next_11,
	out_real_3,
	stg_imag_next_21,
	out_imag_4,
	stg_real_next_21,
	out_real_4,
	stg_imag_next_31,
	out_imag_5,
	stg_real_next_31,
	out_real_5,
	stg_imag_next_41,
	out_imag_6,
	stg_real_next_41,
	out_real_6,
	stg_imag_next_51,
	out_imag_7,
	stg_real_next_51,
	out_real_7,
	stg_imag_next_61,
	out_imag_8,
	stg_real_next_61,
	out_real_8,
	stg_imag_next_71,
	out_imag_9,
	stg_real_next_71,
	out_real_9,
	out_control_2,
	curr_blk_s_1,
	stg_valid_next1,
	out_valid_s,
	out_enable,
	out_valid,
	Equal1,
	stg_inverse_next1,
	out_data_8,
	out_data_0,
	curr_inverse_s,
	out_inverse,
	out_data_9,
	out_data_1,
	out_data_10,
	out_data_2,
	out_data_11,
	out_data_3,
	out_data_12,
	out_data_4,
	out_data_13,
	out_data_5,
	out_data_14,
	out_data_6,
	out_data_15,
	out_data_7,
	stg_in_sop_0,
	out_eop,
	stg_sop_next1,
	stg_eop_next1,
	out_sop,
	out_control_1,
	stg_control_next_1,
	stg_control_next_2,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	stg_imag_next_0;
output 	stg_real_next_0;
output 	stg_imag_next_1;
output 	stg_real_next_1;
output 	stg_imag_next_2;
output 	stg_real_next_2;
output 	stg_imag_next_3;
output 	stg_real_next_3;
output 	stg_imag_next_4;
output 	stg_real_next_4;
output 	stg_imag_next_5;
output 	stg_real_next_5;
output 	stg_imag_next_6;
output 	stg_real_next_6;
output 	stg_imag_next_7;
output 	stg_real_next_7;
output 	stg_imag_next_01;
input 	out_imag_2;
output 	stg_real_next_01;
input 	out_real_2;
output 	stg_imag_next_11;
input 	out_imag_3;
output 	stg_real_next_11;
input 	out_real_3;
output 	stg_imag_next_21;
input 	out_imag_4;
output 	stg_real_next_21;
input 	out_real_4;
output 	stg_imag_next_31;
input 	out_imag_5;
output 	stg_real_next_31;
input 	out_real_5;
output 	stg_imag_next_41;
input 	out_imag_6;
output 	stg_real_next_41;
input 	out_real_6;
output 	stg_imag_next_51;
input 	out_imag_7;
output 	stg_real_next_51;
input 	out_real_7;
output 	stg_imag_next_61;
input 	out_imag_8;
output 	stg_real_next_61;
input 	out_real_8;
output 	stg_imag_next_71;
input 	out_imag_9;
output 	stg_real_next_71;
input 	out_real_9;
input 	out_control_2;
input 	curr_blk_s_1;
output 	stg_valid_next1;
input 	out_valid_s;
input 	out_enable;
input 	out_valid;
input 	Equal1;
output 	stg_inverse_next1;
input 	out_data_8;
input 	out_data_0;
input 	curr_inverse_s;
input 	out_inverse;
input 	out_data_9;
input 	out_data_1;
input 	out_data_10;
input 	out_data_2;
input 	out_data_11;
input 	out_data_3;
input 	out_data_12;
input 	out_data_4;
input 	out_data_13;
input 	out_data_5;
input 	out_data_14;
input 	out_data_6;
input 	out_data_15;
input 	out_data_7;
input 	stg_in_sop_0;
input 	out_eop;
output 	stg_sop_next1;
output 	stg_eop_next1;
input 	out_sop;
input 	out_control_1;
output 	stg_control_next_1;
output 	stg_control_next_2;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \stg_valid_next~0_combout ;
wire \stg_inverse_next~0_combout ;
wire \stg_sop_next~0_combout ;
wire \stg_eop_next~0_combout ;
wire \stg_control_next~0_combout ;
wire \stg_control_next~1_combout ;


dffeas \stg_imag_next[0] (
	.clk(clk),
	.d(stg_imag_next_01),
	.asdata(out_imag_2),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_0),
	.prn(vcc));
defparam \stg_imag_next[0] .is_wysiwyg = "true";
defparam \stg_imag_next[0] .power_up = "low";

dffeas \stg_real_next[0] (
	.clk(clk),
	.d(stg_real_next_01),
	.asdata(out_real_2),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_0),
	.prn(vcc));
defparam \stg_real_next[0] .is_wysiwyg = "true";
defparam \stg_real_next[0] .power_up = "low";

dffeas \stg_imag_next[1] (
	.clk(clk),
	.d(stg_imag_next_11),
	.asdata(out_imag_3),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_1),
	.prn(vcc));
defparam \stg_imag_next[1] .is_wysiwyg = "true";
defparam \stg_imag_next[1] .power_up = "low";

dffeas \stg_real_next[1] (
	.clk(clk),
	.d(stg_real_next_11),
	.asdata(out_real_3),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_1),
	.prn(vcc));
defparam \stg_real_next[1] .is_wysiwyg = "true";
defparam \stg_real_next[1] .power_up = "low";

dffeas \stg_imag_next[2] (
	.clk(clk),
	.d(stg_imag_next_21),
	.asdata(out_imag_4),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_2),
	.prn(vcc));
defparam \stg_imag_next[2] .is_wysiwyg = "true";
defparam \stg_imag_next[2] .power_up = "low";

dffeas \stg_real_next[2] (
	.clk(clk),
	.d(stg_real_next_21),
	.asdata(out_real_4),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_2),
	.prn(vcc));
defparam \stg_real_next[2] .is_wysiwyg = "true";
defparam \stg_real_next[2] .power_up = "low";

dffeas \stg_imag_next[3] (
	.clk(clk),
	.d(stg_imag_next_31),
	.asdata(out_imag_5),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_3),
	.prn(vcc));
defparam \stg_imag_next[3] .is_wysiwyg = "true";
defparam \stg_imag_next[3] .power_up = "low";

dffeas \stg_real_next[3] (
	.clk(clk),
	.d(stg_real_next_31),
	.asdata(out_real_5),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_3),
	.prn(vcc));
defparam \stg_real_next[3] .is_wysiwyg = "true";
defparam \stg_real_next[3] .power_up = "low";

dffeas \stg_imag_next[4] (
	.clk(clk),
	.d(stg_imag_next_41),
	.asdata(out_imag_6),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_4),
	.prn(vcc));
defparam \stg_imag_next[4] .is_wysiwyg = "true";
defparam \stg_imag_next[4] .power_up = "low";

dffeas \stg_real_next[4] (
	.clk(clk),
	.d(stg_real_next_41),
	.asdata(out_real_6),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_4),
	.prn(vcc));
defparam \stg_real_next[4] .is_wysiwyg = "true";
defparam \stg_real_next[4] .power_up = "low";

dffeas \stg_imag_next[5] (
	.clk(clk),
	.d(stg_imag_next_51),
	.asdata(out_imag_7),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_5),
	.prn(vcc));
defparam \stg_imag_next[5] .is_wysiwyg = "true";
defparam \stg_imag_next[5] .power_up = "low";

dffeas \stg_real_next[5] (
	.clk(clk),
	.d(stg_real_next_51),
	.asdata(out_real_7),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_5),
	.prn(vcc));
defparam \stg_real_next[5] .is_wysiwyg = "true";
defparam \stg_real_next[5] .power_up = "low";

dffeas \stg_imag_next[6] (
	.clk(clk),
	.d(stg_imag_next_61),
	.asdata(out_imag_8),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_6),
	.prn(vcc));
defparam \stg_imag_next[6] .is_wysiwyg = "true";
defparam \stg_imag_next[6] .power_up = "low";

dffeas \stg_real_next[6] (
	.clk(clk),
	.d(stg_real_next_61),
	.asdata(out_real_8),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_6),
	.prn(vcc));
defparam \stg_real_next[6] .is_wysiwyg = "true";
defparam \stg_real_next[6] .power_up = "low";

dffeas \stg_imag_next[7] (
	.clk(clk),
	.d(stg_imag_next_71),
	.asdata(out_imag_9),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_imag_next_7),
	.prn(vcc));
defparam \stg_imag_next[7] .is_wysiwyg = "true";
defparam \stg_imag_next[7] .power_up = "low";

dffeas \stg_real_next[7] (
	.clk(clk),
	.d(stg_real_next_71),
	.asdata(out_real_9),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(!curr_blk_s_1),
	.ena(out_enable),
	.q(stg_real_next_7),
	.prn(vcc));
defparam \stg_real_next[7] .is_wysiwyg = "true";
defparam \stg_real_next[7] .power_up = "low";

cycloneiv_lcell_comb \stg_imag_next[0]~0 (
	.dataa(out_data_8),
	.datab(out_data_0),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_01),
	.cout());
defparam \stg_imag_next[0]~0 .lut_mask = 16'hAACC;
defparam \stg_imag_next[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[0]~0 (
	.dataa(out_data_0),
	.datab(out_data_8),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_01),
	.cout());
defparam \stg_real_next[0]~0 .lut_mask = 16'hAACC;
defparam \stg_real_next[0]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[1]~1 (
	.dataa(out_data_9),
	.datab(out_data_1),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_11),
	.cout());
defparam \stg_imag_next[1]~1 .lut_mask = 16'hAACC;
defparam \stg_imag_next[1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[1]~1 (
	.dataa(out_data_1),
	.datab(out_data_9),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_11),
	.cout());
defparam \stg_real_next[1]~1 .lut_mask = 16'hAACC;
defparam \stg_real_next[1]~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[2]~2 (
	.dataa(out_data_10),
	.datab(out_data_2),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_21),
	.cout());
defparam \stg_imag_next[2]~2 .lut_mask = 16'hAACC;
defparam \stg_imag_next[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[2]~2 (
	.dataa(out_data_2),
	.datab(out_data_10),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_21),
	.cout());
defparam \stg_real_next[2]~2 .lut_mask = 16'hAACC;
defparam \stg_real_next[2]~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[3]~3 (
	.dataa(out_data_11),
	.datab(out_data_3),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_31),
	.cout());
defparam \stg_imag_next[3]~3 .lut_mask = 16'hAACC;
defparam \stg_imag_next[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[3]~3 (
	.dataa(out_data_3),
	.datab(out_data_11),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_31),
	.cout());
defparam \stg_real_next[3]~3 .lut_mask = 16'hAACC;
defparam \stg_real_next[3]~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[4]~4 (
	.dataa(out_data_12),
	.datab(out_data_4),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_41),
	.cout());
defparam \stg_imag_next[4]~4 .lut_mask = 16'hAACC;
defparam \stg_imag_next[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[4]~4 (
	.dataa(out_data_4),
	.datab(out_data_12),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_41),
	.cout());
defparam \stg_real_next[4]~4 .lut_mask = 16'hAACC;
defparam \stg_real_next[4]~4 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[5]~5 (
	.dataa(out_data_13),
	.datab(out_data_5),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_51),
	.cout());
defparam \stg_imag_next[5]~5 .lut_mask = 16'hAACC;
defparam \stg_imag_next[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[5]~5 (
	.dataa(out_data_5),
	.datab(out_data_13),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_51),
	.cout());
defparam \stg_real_next[5]~5 .lut_mask = 16'hAACC;
defparam \stg_real_next[5]~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[6]~6 (
	.dataa(out_data_14),
	.datab(out_data_6),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_61),
	.cout());
defparam \stg_imag_next[6]~6 .lut_mask = 16'hAACC;
defparam \stg_imag_next[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[6]~6 (
	.dataa(out_data_6),
	.datab(out_data_14),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_61),
	.cout());
defparam \stg_real_next[6]~6 .lut_mask = 16'hAACC;
defparam \stg_real_next[6]~6 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_imag_next[7]~7 (
	.dataa(out_data_15),
	.datab(out_data_7),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_imag_next_71),
	.cout());
defparam \stg_imag_next[7]~7 .lut_mask = 16'hAACC;
defparam \stg_imag_next[7]~7 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_real_next[7]~7 (
	.dataa(out_data_7),
	.datab(out_data_15),
	.datac(gnd),
	.datad(curr_inverse_s),
	.cin(gnd),
	.combout(stg_real_next_71),
	.cout());
defparam \stg_real_next[7]~7 .lut_mask = 16'hAACC;
defparam \stg_real_next[7]~7 .sum_lutc_input = "datac";

dffeas stg_valid_next(
	.clk(clk),
	.d(\stg_valid_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_valid_next1),
	.prn(vcc));
defparam stg_valid_next.is_wysiwyg = "true";
defparam stg_valid_next.power_up = "low";

dffeas stg_inverse_next(
	.clk(clk),
	.d(\stg_inverse_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_inverse_next1),
	.prn(vcc));
defparam stg_inverse_next.is_wysiwyg = "true";
defparam stg_inverse_next.power_up = "low";

dffeas stg_sop_next(
	.clk(clk),
	.d(\stg_sop_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_sop_next1),
	.prn(vcc));
defparam stg_sop_next.is_wysiwyg = "true";
defparam stg_sop_next.power_up = "low";

dffeas stg_eop_next(
	.clk(clk),
	.d(\stg_eop_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_eop_next1),
	.prn(vcc));
defparam stg_eop_next.is_wysiwyg = "true";
defparam stg_eop_next.power_up = "low";

dffeas \stg_control_next[1] (
	.clk(clk),
	.d(\stg_control_next~0_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_control_next_1),
	.prn(vcc));
defparam \stg_control_next[1] .is_wysiwyg = "true";
defparam \stg_control_next[1] .power_up = "low";

dffeas \stg_control_next[2] (
	.clk(clk),
	.d(\stg_control_next~1_combout ),
	.asdata(vcc),
	.clrn(reset_n),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(out_enable),
	.q(stg_control_next_2),
	.prn(vcc));
defparam \stg_control_next[2] .is_wysiwyg = "true";
defparam \stg_control_next[2] .power_up = "low";

cycloneiv_lcell_comb \stg_valid_next~0 (
	.dataa(out_valid_s),
	.datab(out_valid),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_valid_next~0_combout ),
	.cout());
defparam \stg_valid_next~0 .lut_mask = 16'hAACC;
defparam \stg_valid_next~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_inverse_next~0 (
	.dataa(curr_inverse_s),
	.datab(out_inverse),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_inverse_next~0_combout ),
	.cout());
defparam \stg_inverse_next~0 .lut_mask = 16'hAACC;
defparam \stg_inverse_next~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_sop_next~0 (
	.dataa(stg_in_sop_0),
	.datab(out_sop),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_sop_next~0_combout ),
	.cout());
defparam \stg_sop_next~0 .lut_mask = 16'hAACC;
defparam \stg_sop_next~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_eop_next~0 (
	.dataa(Equal1),
	.datab(out_eop),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_eop_next~0_combout ),
	.cout());
defparam \stg_eop_next~0 .lut_mask = 16'hCC55;
defparam \stg_eop_next~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_control_next~0 (
	.dataa(out_control_1),
	.datab(gnd),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_control_next~0_combout ),
	.cout());
defparam \stg_control_next~0 .lut_mask = 16'hAAFF;
defparam \stg_control_next~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \stg_control_next~1 (
	.dataa(out_control_2),
	.datab(gnd),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\stg_control_next~1_combout ),
	.cout());
defparam \stg_control_next~1 .lut_mask = 16'hAAFF;
defparam \stg_control_next~1 .sum_lutc_input = "datac";

endmodule

module ifft_8p_auk_dspip_r22sdf_twrom (
	imagtwid_0,
	imagtwid_1,
	imagtwid_2,
	imagtwid_3,
	imagtwid_4,
	imagtwid_5,
	imagtwid_6,
	imagtwid_7,
	curr_blk_s_1,
	stg_valid_next,
	curr_pwr_2_s,
	enable,
	realtwid_0,
	realtwid_1,
	realtwid_2,
	realtwid_3,
	realtwid_4,
	realtwid_5,
	realtwid_6,
	realtwid_7,
	control_s_1,
	control_s_2,
	control_s_0,
	rd_en,
	GND_port,
	clk,
	reset)/* synthesis synthesis_greybox=1 */;
output 	imagtwid_0;
output 	imagtwid_1;
output 	imagtwid_2;
output 	imagtwid_3;
output 	imagtwid_4;
output 	imagtwid_5;
output 	imagtwid_6;
output 	imagtwid_7;
input 	curr_blk_s_1;
input 	stg_valid_next;
input 	curr_pwr_2_s;
input 	enable;
output 	realtwid_0;
output 	realtwid_1;
output 	realtwid_2;
output 	realtwid_3;
output 	realtwid_4;
output 	realtwid_5;
output 	realtwid_6;
output 	realtwid_7;
input 	control_s_1;
input 	control_s_2;
input 	control_s_0;
input 	rd_en;
input 	GND_port;
input 	clk;
input 	reset;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;

wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ;
wire \gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ;
wire \gen_optimized_memory_delayed:addr_real_s[1]~0_combout ;
wire \gen_optimized_memory_delayed:addr_imag_s[1]~0_combout ;
wire \imagtwid[0]~8_combout ;
wire \cnt_grp~0_combout ;
wire \gen_optimized_memory_delayed:cnt_grp[1]~0_combout ;
wire \gen_optimized_memory_delayed:cnt_grp_d[0][1]~q ;
wire \gen_optimized_memory_delayed:cnt_grp_d[1][1]~q ;
wire \gen_optimized_memory_delayed:cnt_grp[0]~0_combout ;
wire \gen_optimized_memory_delayed:cnt_grp_d[0][0]~q ;
wire \gen_optimized_memory_delayed:cnt_grp_d[1][0]~q ;
wire \Equal1~0_combout ;
wire \Mux0~0_combout ;
wire \gen_optimized_memory_delayed:cnt_w_k[0]~1_combout ;
wire \gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d~q ;
wire \cnt_w_k~0_combout ;
wire \cnt_w_k~1_combout ;
wire \cnt_w_k~2_combout ;
wire \cnt_w_k~3_combout ;
wire \cnt_w_k~4_combout ;
wire \gen_optimized_memory_delayed:cnt_w_k[0]~q ;
wire \gen_optimized_memory_delayed:cnt_w_k[0]~2 ;
wire \gen_optimized_memory_delayed:cnt_w_k[1]~1_combout ;
wire \Add1~0_combout ;
wire \gen_optimized_memory_delayed:cnt_w_k[1]~q ;
wire \gen_optimized_memory_delayed:cnt_w_k[1]~2 ;
wire \gen_optimized_memory_delayed:cnt_w_k[2]~1_combout ;
wire \Add1~1_combout ;
wire \gen_optimized_memory_delayed:cnt_w_k[2]~q ;
wire \gen_optimized_memory_delayed:negate_op_d[0][1]~q ;
wire \gen_optimized_memory_delayed:negate_op_d[1][1]~q ;
wire \imagtwid[0]~9 ;
wire \imagtwid[1]~10_combout ;
wire \imagtwid[1]~11 ;
wire \imagtwid[2]~12_combout ;
wire \imagtwid[2]~13 ;
wire \imagtwid[3]~14_combout ;
wire \imagtwid[3]~15 ;
wire \imagtwid[4]~16_combout ;
wire \imagtwid[4]~17 ;
wire \imagtwid[5]~18_combout ;
wire \imagtwid[5]~19 ;
wire \imagtwid[6]~20_combout ;
wire \imagtwid[6]~21 ;
wire \imagtwid[0]~23_cout ;
wire \imagtwid[7]~24_combout ;
wire \Add4~0_combout ;
wire \Add4~2_cout ;
wire \Add4~3_combout ;
wire \gen_optimized_memory_delayed:negate_op_d[0][0]~q ;
wire \gen_optimized_memory_delayed:negate_op_d[1][0]~q ;
wire \reg_negate_op~0_combout ;
wire \Add4~5_combout ;
wire \Add4~4 ;
wire \Add4~6_combout ;
wire \Add4~8_combout ;
wire \Add4~7 ;
wire \Add4~9_combout ;
wire \Add4~11_combout ;
wire \Add4~10 ;
wire \Add4~12_combout ;
wire \Add4~14_combout ;
wire \Add4~13 ;
wire \Add4~15_combout ;
wire \Add4~17_combout ;
wire \Add4~16 ;
wire \Add4~18_combout ;
wire \Add4~20_combout ;
wire \Add4~19 ;
wire \Add4~22_cout ;
wire \Add4~23_combout ;
wire \Add4~25_combout ;


ifft_8p_altera_fft_dual_port_rom \gen_optimized_memory_delayed:dual_port_rom_component (
	.q_a_0(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.q_b_0(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.q_a_1(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.q_b_1(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.q_a_2(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.q_b_2(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.q_a_3(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.q_b_3(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.q_a_4(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.q_b_4(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.q_a_5(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.q_b_5(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.q_a_6(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.q_b_6(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.q_a_7(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.q_b_7(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.gen_optimized_memory_delayedcnt_w_k0(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.out_enable(enable),
	.gen_optimized_memory_delayedaddr_real_s1(\gen_optimized_memory_delayed:addr_real_s[1]~0_combout ),
	.gen_optimized_memory_delayedaddr_imag_s1(\gen_optimized_memory_delayed:addr_imag_s[1]~0_combout ),
	.GND_port(GND_port),
	.clk(clk),
	.reset_n(reset));

cycloneiv_lcell_comb \gen_optimized_memory_delayed:addr_real_s[1]~0 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.cin(gnd),
	.combout(\gen_optimized_memory_delayed:addr_real_s[1]~0_combout ),
	.cout());
defparam \gen_optimized_memory_delayed:addr_real_s[1]~0 .lut_mask = 16'hFF55;
defparam \gen_optimized_memory_delayed:addr_real_s[1]~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:addr_imag_s[1]~0 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.datab(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\gen_optimized_memory_delayed:addr_imag_s[1]~0_combout ),
	.cout());
defparam \gen_optimized_memory_delayed:addr_imag_s[1]~0 .lut_mask = 16'h7777;
defparam \gen_optimized_memory_delayed:addr_imag_s[1]~0 .sum_lutc_input = "datac";

dffeas \imagtwid[0] (
	.clk(clk),
	.d(\imagtwid[0]~8_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_0),
	.prn(vcc));
defparam \imagtwid[0] .is_wysiwyg = "true";
defparam \imagtwid[0] .power_up = "low";

dffeas \imagtwid[1] (
	.clk(clk),
	.d(\imagtwid[1]~10_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_1),
	.prn(vcc));
defparam \imagtwid[1] .is_wysiwyg = "true";
defparam \imagtwid[1] .power_up = "low";

dffeas \imagtwid[2] (
	.clk(clk),
	.d(\imagtwid[2]~12_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_2),
	.prn(vcc));
defparam \imagtwid[2] .is_wysiwyg = "true";
defparam \imagtwid[2] .power_up = "low";

dffeas \imagtwid[3] (
	.clk(clk),
	.d(\imagtwid[3]~14_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_3),
	.prn(vcc));
defparam \imagtwid[3] .is_wysiwyg = "true";
defparam \imagtwid[3] .power_up = "low";

dffeas \imagtwid[4] (
	.clk(clk),
	.d(\imagtwid[4]~16_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_4),
	.prn(vcc));
defparam \imagtwid[4] .is_wysiwyg = "true";
defparam \imagtwid[4] .power_up = "low";

dffeas \imagtwid[5] (
	.clk(clk),
	.d(\imagtwid[5]~18_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_5),
	.prn(vcc));
defparam \imagtwid[5] .is_wysiwyg = "true";
defparam \imagtwid[5] .power_up = "low";

dffeas \imagtwid[6] (
	.clk(clk),
	.d(\imagtwid[6]~20_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_6),
	.prn(vcc));
defparam \imagtwid[6] .is_wysiwyg = "true";
defparam \imagtwid[6] .power_up = "low";

dffeas \imagtwid[7] (
	.clk(clk),
	.d(\imagtwid[7]~24_combout ),
	.asdata(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\Equal1~0_combout ),
	.sload(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.ena(enable),
	.q(imagtwid_7),
	.prn(vcc));
defparam \imagtwid[7] .is_wysiwyg = "true";
defparam \imagtwid[7] .power_up = "low";

dffeas \realtwid[0] (
	.clk(clk),
	.d(\Add4~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_0),
	.prn(vcc));
defparam \realtwid[0] .is_wysiwyg = "true";
defparam \realtwid[0] .power_up = "low";

dffeas \realtwid[1] (
	.clk(clk),
	.d(\Add4~5_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_1),
	.prn(vcc));
defparam \realtwid[1] .is_wysiwyg = "true";
defparam \realtwid[1] .power_up = "low";

dffeas \realtwid[2] (
	.clk(clk),
	.d(\Add4~8_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_2),
	.prn(vcc));
defparam \realtwid[2] .is_wysiwyg = "true";
defparam \realtwid[2] .power_up = "low";

dffeas \realtwid[3] (
	.clk(clk),
	.d(\Add4~11_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_3),
	.prn(vcc));
defparam \realtwid[3] .is_wysiwyg = "true";
defparam \realtwid[3] .power_up = "low";

dffeas \realtwid[4] (
	.clk(clk),
	.d(\Add4~14_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_4),
	.prn(vcc));
defparam \realtwid[4] .is_wysiwyg = "true";
defparam \realtwid[4] .power_up = "low";

dffeas \realtwid[5] (
	.clk(clk),
	.d(\Add4~17_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_5),
	.prn(vcc));
defparam \realtwid[5] .is_wysiwyg = "true";
defparam \realtwid[5] .power_up = "low";

dffeas \realtwid[6] (
	.clk(clk),
	.d(\Add4~20_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_6),
	.prn(vcc));
defparam \realtwid[6] .is_wysiwyg = "true";
defparam \realtwid[6] .power_up = "low";

dffeas \realtwid[7] (
	.clk(clk),
	.d(\Add4~25_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(realtwid_7),
	.prn(vcc));
defparam \realtwid[7] .is_wysiwyg = "true";
defparam \realtwid[7] .power_up = "low";

cycloneiv_lcell_comb \imagtwid[0]~8 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\imagtwid[0]~8_combout ),
	.cout(\imagtwid[0]~9 ));
defparam \imagtwid[0]~8 .lut_mask = 16'hAA55;
defparam \imagtwid[0]~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt_grp~0 (
	.dataa(curr_blk_s_1),
	.datab(curr_pwr_2_s),
	.datac(stg_valid_next),
	.datad(control_s_0),
	.cin(gnd),
	.combout(\cnt_grp~0_combout ),
	.cout());
defparam \cnt_grp~0 .lut_mask = 16'hBFFF;
defparam \cnt_grp~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:cnt_grp[1]~0 (
	.dataa(\cnt_grp~0_combout ),
	.datab(control_s_2),
	.datac(control_s_1),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\gen_optimized_memory_delayed:cnt_grp[1]~0_combout ),
	.cout());
defparam \gen_optimized_memory_delayed:cnt_grp[1]~0 .lut_mask = 16'hAFCF;
defparam \gen_optimized_memory_delayed:cnt_grp[1]~0 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:cnt_grp_d[0][1] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_grp[1]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_grp_d[0][1]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_grp_d[0][1] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_grp_d[0][1] .power_up = "low";

dffeas \gen_optimized_memory_delayed:cnt_grp_d[1][1] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_grp_d[0][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_grp_d[1][1]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_grp_d[1][1] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_grp_d[1][1] .power_up = "low";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:cnt_grp[0]~0 (
	.dataa(\cnt_grp~0_combout ),
	.datab(control_s_1),
	.datac(control_s_2),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\gen_optimized_memory_delayed:cnt_grp[0]~0_combout ),
	.cout());
defparam \gen_optimized_memory_delayed:cnt_grp[0]~0 .lut_mask = 16'hAFCF;
defparam \gen_optimized_memory_delayed:cnt_grp[0]~0 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:cnt_grp_d[0][0] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_grp[0]~0_combout ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_grp_d[0][0]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_grp_d[0][0] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_grp_d[0][0] .power_up = "low";

dffeas \gen_optimized_memory_delayed:cnt_grp_d[1][0] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_grp_d[0][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_grp_d[1][0]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_grp_d[1][0] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_grp_d[1][0] .power_up = "low";

cycloneiv_lcell_comb \Equal1~0 (
	.dataa(\gen_optimized_memory_delayed:cnt_grp_d[1][1]~q ),
	.datab(\gen_optimized_memory_delayed:cnt_grp_d[1][0]~q ),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
defparam \Equal1~0 .lut_mask = 16'hEEEE;
defparam \Equal1~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Mux0~0 (
	.dataa(control_s_1),
	.datab(control_s_2),
	.datac(curr_blk_s_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
defparam \Mux0~0 .lut_mask = 16'h6F6F;
defparam \Mux0~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:cnt_w_k[0]~1 (
	.dataa(\Mux0~0_combout ),
	.datab(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\gen_optimized_memory_delayed:cnt_w_k[0]~1_combout ),
	.cout(\gen_optimized_memory_delayed:cnt_w_k[0]~2 ));
defparam \gen_optimized_memory_delayed:cnt_w_k[0]~1 .lut_mask = 16'h66EE;
defparam \gen_optimized_memory_delayed:cnt_w_k[0]~1 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d (
	.clk(clk),
	.d(rd_en),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d .power_up = "low";

cycloneiv_lcell_comb \cnt_w_k~0 (
	.dataa(\gen_optimized_memory_delayed:gen_max_pwr_2:rd_en_d~q ),
	.datab(curr_pwr_2_s),
	.datac(curr_blk_s_1),
	.datad(control_s_0),
	.cin(gnd),
	.combout(\cnt_w_k~0_combout ),
	.cout());
defparam \cnt_w_k~0 .lut_mask = 16'hEBBE;
defparam \cnt_w_k~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt_w_k~1 (
	.dataa(control_s_2),
	.datab(control_s_1),
	.datac(gnd),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\cnt_w_k~1_combout ),
	.cout());
defparam \cnt_w_k~1 .lut_mask = 16'hBBFF;
defparam \cnt_w_k~1 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt_w_k~2 (
	.dataa(control_s_2),
	.datab(control_s_1),
	.datac(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\cnt_w_k~2_combout ),
	.cout());
defparam \cnt_w_k~2 .lut_mask = 16'h96FF;
defparam \cnt_w_k~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt_w_k~3 (
	.dataa(\gen_optimized_memory_delayed:cnt_grp[1]~0_combout ),
	.datab(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.datac(\cnt_w_k~1_combout ),
	.datad(\cnt_w_k~2_combout ),
	.cin(gnd),
	.combout(\cnt_w_k~3_combout ),
	.cout());
defparam \cnt_w_k~3 .lut_mask = 16'hEBBE;
defparam \cnt_w_k~3 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \cnt_w_k~4 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[2]~q ),
	.datab(\cnt_w_k~0_combout ),
	.datac(\cnt_w_k~1_combout ),
	.datad(\cnt_w_k~3_combout ),
	.cin(gnd),
	.combout(\cnt_w_k~4_combout ),
	.cout());
defparam \cnt_w_k~4 .lut_mask = 16'hFBFF;
defparam \cnt_w_k~4 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:cnt_w_k[0] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_w_k[0]~1_combout ),
	.asdata(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\cnt_w_k~4_combout ),
	.sload(!curr_pwr_2_s),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_w_k[0]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_w_k[0] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_w_k[0] .power_up = "low";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:cnt_w_k[1]~1 (
	.dataa(\gen_optimized_memory_delayed:cnt_grp[0]~0_combout ),
	.datab(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.datac(gnd),
	.datad(vcc),
	.cin(\gen_optimized_memory_delayed:cnt_w_k[0]~2 ),
	.combout(\gen_optimized_memory_delayed:cnt_w_k[1]~1_combout ),
	.cout(\gen_optimized_memory_delayed:cnt_w_k[1]~2 ));
defparam \gen_optimized_memory_delayed:cnt_w_k[1]~1 .lut_mask = 16'h96BF;
defparam \gen_optimized_memory_delayed:cnt_w_k[1]~1 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add1~0 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.datab(control_s_1),
	.datac(control_s_2),
	.datad(curr_blk_s_1),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout());
defparam \Add1~0 .lut_mask = 16'h6996;
defparam \Add1~0 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:cnt_w_k[1] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_w_k[1]~1_combout ),
	.asdata(\Add1~0_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\cnt_w_k~4_combout ),
	.sload(!curr_pwr_2_s),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_w_k[1] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_w_k[1] .power_up = "low";

cycloneiv_lcell_comb \gen_optimized_memory_delayed:cnt_w_k[2]~1 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[2]~q ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\gen_optimized_memory_delayed:cnt_w_k[1]~2 ),
	.combout(\gen_optimized_memory_delayed:cnt_w_k[2]~1_combout ),
	.cout());
defparam \gen_optimized_memory_delayed:cnt_w_k[2]~1 .lut_mask = 16'h5A5A;
defparam \gen_optimized_memory_delayed:cnt_w_k[2]~1 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add1~1 (
	.dataa(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.datab(\Mux0~0_combout ),
	.datac(\gen_optimized_memory_delayed:cnt_grp[0]~0_combout ),
	.datad(\gen_optimized_memory_delayed:cnt_w_k[2]~q ),
	.cin(gnd),
	.combout(\Add1~1_combout ),
	.cout());
defparam \Add1~1 .lut_mask = 16'h6996;
defparam \Add1~1 .sum_lutc_input = "datac";

dffeas \gen_optimized_memory_delayed:cnt_w_k[2] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_w_k[2]~1_combout ),
	.asdata(\Add1~1_combout ),
	.clrn(reset),
	.aload(gnd),
	.sclr(\cnt_w_k~4_combout ),
	.sload(!curr_pwr_2_s),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:cnt_w_k[2]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:cnt_w_k[2] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:cnt_w_k[2] .power_up = "low";

dffeas \gen_optimized_memory_delayed:negate_op_d[0][1] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_w_k[2]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:negate_op_d[0][1]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:negate_op_d[0][1] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:negate_op_d[0][1] .power_up = "low";

dffeas \gen_optimized_memory_delayed:negate_op_d[1][1] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:negate_op_d[0][1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:negate_op_d[1][1] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:negate_op_d[1][1] .power_up = "low";

cycloneiv_lcell_comb \imagtwid[1]~10 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[0]~9 ),
	.combout(\imagtwid[1]~10_combout ),
	.cout(\imagtwid[1]~11 ));
defparam \imagtwid[1]~10 .lut_mask = 16'h5AAF;
defparam \imagtwid[1]~10 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[2]~12 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[1]~11 ),
	.combout(\imagtwid[2]~12_combout ),
	.cout(\imagtwid[2]~13 ));
defparam \imagtwid[2]~12 .lut_mask = 16'h5A5F;
defparam \imagtwid[2]~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[3]~14 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[2]~13 ),
	.combout(\imagtwid[3]~14_combout ),
	.cout(\imagtwid[3]~15 ));
defparam \imagtwid[3]~14 .lut_mask = 16'h5AAF;
defparam \imagtwid[3]~14 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[4]~16 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[3]~15 ),
	.combout(\imagtwid[4]~16_combout ),
	.cout(\imagtwid[4]~17 ));
defparam \imagtwid[4]~16 .lut_mask = 16'h5A5F;
defparam \imagtwid[4]~16 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[5]~18 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[4]~17 ),
	.combout(\imagtwid[5]~18_combout ),
	.cout(\imagtwid[5]~19 ));
defparam \imagtwid[5]~18 .lut_mask = 16'h5AAF;
defparam \imagtwid[5]~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[6]~20 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[5]~19 ),
	.combout(\imagtwid[6]~20_combout ),
	.cout(\imagtwid[6]~21 ));
defparam \imagtwid[6]~20 .lut_mask = 16'h5A5F;
defparam \imagtwid[6]~20 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[0]~23 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\imagtwid[6]~21 ),
	.combout(),
	.cout(\imagtwid[0]~23_cout ));
defparam \imagtwid[0]~23 .lut_mask = 16'h00AF;
defparam \imagtwid[0]~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \imagtwid[7]~24 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_b[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\imagtwid[0]~23_cout ),
	.combout(\imagtwid[7]~24_combout ),
	.cout());
defparam \imagtwid[7]~24 .lut_mask = 16'h5A5A;
defparam \imagtwid[7]~24 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~0 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datab(\gen_optimized_memory_delayed:cnt_grp_d[1][1]~q ),
	.datac(\gen_optimized_memory_delayed:cnt_grp_d[1][0]~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\Add4~0_combout ),
	.cout());
defparam \Add4~0 .lut_mask = 16'hFEFE;
defparam \Add4~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~2 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[0] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\Add4~2_cout ));
defparam \Add4~2 .lut_mask = 16'h0055;
defparam \Add4~2 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~3 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~2_cout ),
	.combout(\Add4~3_combout ),
	.cout(\Add4~4 ));
defparam \Add4~3 .lut_mask = 16'h5AAF;
defparam \Add4~3 .sum_lutc_input = "cin";

dffeas \gen_optimized_memory_delayed:negate_op_d[0][0] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:cnt_w_k[1]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:negate_op_d[0][0]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:negate_op_d[0][0] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:negate_op_d[0][0] .power_up = "low";

dffeas \gen_optimized_memory_delayed:negate_op_d[1][0] (
	.clk(clk),
	.d(\gen_optimized_memory_delayed:negate_op_d[0][0]~q ),
	.asdata(vcc),
	.clrn(reset),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(enable),
	.q(\gen_optimized_memory_delayed:negate_op_d[1][0]~q ),
	.prn(vcc));
defparam \gen_optimized_memory_delayed:negate_op_d[1][0] .is_wysiwyg = "true";
defparam \gen_optimized_memory_delayed:negate_op_d[1][0] .power_up = "low";

cycloneiv_lcell_comb \reg_negate_op~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\gen_optimized_memory_delayed:negate_op_d[1][1]~q ),
	.datad(\gen_optimized_memory_delayed:negate_op_d[1][0]~q ),
	.cin(gnd),
	.combout(\reg_negate_op~0_combout ),
	.cout());
defparam \reg_negate_op~0 .lut_mask = 16'h0FF0;
defparam \reg_negate_op~0 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~5 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~3_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[1] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~5_combout ),
	.cout());
defparam \Add4~5 .lut_mask = 16'hFAFC;
defparam \Add4~5 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~6 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~4 ),
	.combout(\Add4~6_combout ),
	.cout(\Add4~7 ));
defparam \Add4~6 .lut_mask = 16'h5A5F;
defparam \Add4~6 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~8 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~6_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[2] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~8_combout ),
	.cout());
defparam \Add4~8 .lut_mask = 16'hFAFC;
defparam \Add4~8 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~9 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~7 ),
	.combout(\Add4~9_combout ),
	.cout(\Add4~10 ));
defparam \Add4~9 .lut_mask = 16'h5AAF;
defparam \Add4~9 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~11 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~9_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[3] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~11_combout ),
	.cout());
defparam \Add4~11 .lut_mask = 16'hFAFC;
defparam \Add4~11 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~12 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~10 ),
	.combout(\Add4~12_combout ),
	.cout(\Add4~13 ));
defparam \Add4~12 .lut_mask = 16'h5A5F;
defparam \Add4~12 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~14 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~12_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[4] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~14_combout ),
	.cout());
defparam \Add4~14 .lut_mask = 16'hFAFC;
defparam \Add4~14 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~15 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~13 ),
	.combout(\Add4~15_combout ),
	.cout(\Add4~16 ));
defparam \Add4~15 .lut_mask = 16'h5AAF;
defparam \Add4~15 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~17 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~15_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[5] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~17_combout ),
	.cout());
defparam \Add4~17 .lut_mask = 16'hFAFC;
defparam \Add4~17 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~18 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~16 ),
	.combout(\Add4~18_combout ),
	.cout(\Add4~19 ));
defparam \Add4~18 .lut_mask = 16'h5A5F;
defparam \Add4~18 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~20 (
	.dataa(\Equal1~0_combout ),
	.datab(\Add4~18_combout ),
	.datac(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[6] ),
	.datad(\reg_negate_op~0_combout ),
	.cin(gnd),
	.combout(\Add4~20_combout ),
	.cout());
defparam \Add4~20 .lut_mask = 16'hFAFC;
defparam \Add4~20 .sum_lutc_input = "datac";

cycloneiv_lcell_comb \Add4~22 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add4~19 ),
	.combout(),
	.cout(\Add4~22_cout ));
defparam \Add4~22 .lut_mask = 16'h00AF;
defparam \Add4~22 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~23 (
	.dataa(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add4~22_cout ),
	.combout(\Add4~23_combout ),
	.cout());
defparam \Add4~23 .lut_mask = 16'h5A5A;
defparam \Add4~23 .sum_lutc_input = "cin";

cycloneiv_lcell_comb \Add4~25 (
	.dataa(\Add4~23_combout ),
	.datab(\gen_optimized_memory_delayed:dual_port_rom_component|old_ram_gen:old_ram_component|auto_generated|q_a[7] ),
	.datac(\reg_negate_op~0_combout ),
	.datad(\Equal1~0_combout ),
	.cin(gnd),
	.combout(\Add4~25_combout ),
	.cout());
defparam \Add4~25 .lut_mask = 16'hACFF;
defparam \Add4~25 .sum_lutc_input = "datac";

endmodule

module ifft_8p_altera_fft_dual_port_rom (
	q_a_0,
	q_b_0,
	q_a_1,
	q_b_1,
	q_a_2,
	q_b_2,
	q_a_3,
	q_b_3,
	q_a_4,
	q_b_4,
	q_a_5,
	q_b_5,
	q_a_6,
	q_b_6,
	q_a_7,
	q_b_7,
	gen_optimized_memory_delayedcnt_w_k0,
	out_enable,
	gen_optimized_memory_delayedaddr_real_s1,
	gen_optimized_memory_delayedaddr_imag_s1,
	GND_port,
	clk,
	reset_n)/* synthesis synthesis_greybox=1 */;
output 	q_a_0;
output 	q_b_0;
output 	q_a_1;
output 	q_b_1;
output 	q_a_2;
output 	q_b_2;
output 	q_a_3;
output 	q_b_3;
output 	q_a_4;
output 	q_b_4;
output 	q_a_5;
output 	q_b_5;
output 	q_a_6;
output 	q_b_6;
output 	q_a_7;
output 	q_b_7;
input 	gen_optimized_memory_delayedcnt_w_k0;
input 	out_enable;
input 	gen_optimized_memory_delayedaddr_real_s1;
input 	gen_optimized_memory_delayedaddr_imag_s1;
input 	GND_port;
input 	clk;
input 	reset_n;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altsyncram_2 \old_ram_gen:old_ram_component (
	.q_a({q_a_unconnected_wire_15,q_a_unconnected_wire_14,q_a_unconnected_wire_13,q_a_unconnected_wire_12,q_a_unconnected_wire_11,q_a_unconnected_wire_10,q_a_unconnected_wire_9,q_a_unconnected_wire_8,q_a_7,q_a_6,q_a_5,q_a_4,q_a_3,q_a_2,q_a_1,q_a_0}),
	.q_b({q_b_unconnected_wire_15,q_b_unconnected_wire_14,q_b_unconnected_wire_13,q_b_unconnected_wire_12,q_b_unconnected_wire_11,q_b_unconnected_wire_10,q_b_unconnected_wire_9,q_b_unconnected_wire_8,q_b_7,q_b_6,q_b_5,q_b_4,q_b_3,q_b_2,q_b_1,q_b_0}),
	.address_a({gnd,gen_optimized_memory_delayedaddr_real_s1,gen_optimized_memory_delayedcnt_w_k0}),
	.clocken0(out_enable),
	.address_b({gnd,gen_optimized_memory_delayedaddr_imag_s1,gnd}),
	.data_a({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,GND_port}),
	.clock0(clk),
	.aclr0(reset_n));

endmodule

module ifft_8p_altsyncram_2 (
	q_a,
	q_b,
	address_a,
	clocken0,
	address_b,
	data_a,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	[15:0] q_a;
output 	[15:0] q_b;
input 	[2:0] address_a;
input 	clocken0;
input 	[2:0] address_b;
input 	[15:0] data_a;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;



ifft_8p_altsyncram_obt3 auto_generated(
	.q_a({q_a[7],q_a[6],q_a[5],q_a[4],q_a[3],q_a[2],q_a[1],q_a[0]}),
	.q_b({q_b[7],q_b[6],q_b[5],q_b[4],q_b[3],q_b[2],q_b[1],q_b[0]}),
	.address_a({address_a[1],address_a[0]}),
	.address_b({address_b[1],address_a[0]}),
	.clocken0(clocken0),
	.data_a({data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0]}),
	.data_b({data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0],data_a[0]}),
	.clock0(clock0),
	.aclr0(aclr0));

endmodule

module ifft_8p_altsyncram_obt3 (
	q_a,
	q_b,
	address_a,
	address_b,
	clocken0,
	data_a,
	data_b,
	clock0,
	aclr0)/* synthesis synthesis_greybox=1 */;
output 	[7:0] q_a;
output 	[7:0] q_b;
input 	[1:0] address_a;
input 	[1:0] address_b;
input 	clocken0;
input 	[7:0] data_a;
input 	[7:0] data_b;
input 	clock0;
input 	aclr0;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
// unknown value (1'bx) is not needed for this tool. Default to 1'b0
assign unknown = 1'b0;


wire [143:0] ram_block1a0_PORTADATAOUT_bus;
wire [143:0] ram_block1a0_PORTBDATAOUT_bus;
wire [143:0] ram_block1a1_PORTADATAOUT_bus;
wire [143:0] ram_block1a1_PORTBDATAOUT_bus;
wire [143:0] ram_block1a2_PORTADATAOUT_bus;
wire [143:0] ram_block1a2_PORTBDATAOUT_bus;
wire [143:0] ram_block1a3_PORTADATAOUT_bus;
wire [143:0] ram_block1a3_PORTBDATAOUT_bus;
wire [143:0] ram_block1a4_PORTADATAOUT_bus;
wire [143:0] ram_block1a4_PORTBDATAOUT_bus;
wire [143:0] ram_block1a5_PORTADATAOUT_bus;
wire [143:0] ram_block1a5_PORTBDATAOUT_bus;
wire [143:0] ram_block1a6_PORTADATAOUT_bus;
wire [143:0] ram_block1a6_PORTBDATAOUT_bus;
wire [143:0] ram_block1a7_PORTADATAOUT_bus;
wire [143:0] ram_block1a7_PORTBDATAOUT_bus;

assign q_a[0] = ram_block1a0_PORTADATAOUT_bus[0];

assign q_b[0] = ram_block1a0_PORTBDATAOUT_bus[0];

assign q_a[1] = ram_block1a1_PORTADATAOUT_bus[0];

assign q_b[1] = ram_block1a1_PORTBDATAOUT_bus[0];

assign q_a[2] = ram_block1a2_PORTADATAOUT_bus[0];

assign q_b[2] = ram_block1a2_PORTBDATAOUT_bus[0];

assign q_a[3] = ram_block1a3_PORTADATAOUT_bus[0];

assign q_b[3] = ram_block1a3_PORTBDATAOUT_bus[0];

assign q_a[4] = ram_block1a4_PORTADATAOUT_bus[0];

assign q_b[4] = ram_block1a4_PORTBDATAOUT_bus[0];

assign q_a[5] = ram_block1a5_PORTADATAOUT_bus[0];

assign q_b[5] = ram_block1a5_PORTBDATAOUT_bus[0];

assign q_a[6] = ram_block1a6_PORTADATAOUT_bus[0];

assign q_b[6] = ram_block1a6_PORTBDATAOUT_bus[0];

assign q_a[7] = ram_block1a7_PORTADATAOUT_bus[0];

assign q_b[7] = ram_block1a7_PORTBDATAOUT_bus[0];

cycloneiv_ram_block ram_block1a0(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a0_PORTADATAOUT_bus),
	.portbdataout(ram_block1a0_PORTBDATAOUT_bus));
defparam ram_block1a0.clk0_core_clock_enable = "ena0";
defparam ram_block1a0.clk0_input_clock_enable = "ena0";
defparam ram_block1a0.clk0_output_clock_enable = "ena0";
defparam ram_block1a0.data_interleave_offset_in_bits = 1;
defparam ram_block1a0.data_interleave_width_in_bits = 1;
defparam ram_block1a0.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a0.init_file_layout = "port_a";
defparam ram_block1a0.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a0.operation_mode = "bidir_dual_port";
defparam ram_block1a0.port_a_address_clear = "none";
defparam ram_block1a0.port_a_address_width = 2;
defparam ram_block1a0.port_a_data_out_clear = "clear0";
defparam ram_block1a0.port_a_data_out_clock = "clock0";
defparam ram_block1a0.port_a_data_width = 1;
defparam ram_block1a0.port_a_first_address = 0;
defparam ram_block1a0.port_a_first_bit_number = 0;
defparam ram_block1a0.port_a_last_address = 2;
defparam ram_block1a0.port_a_logical_ram_depth = 3;
defparam ram_block1a0.port_a_logical_ram_width = 8;
defparam ram_block1a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_address_clear = "none";
defparam ram_block1a0.port_b_address_clock = "clock0";
defparam ram_block1a0.port_b_address_width = 2;
defparam ram_block1a0.port_b_data_in_clock = "clock0";
defparam ram_block1a0.port_b_data_out_clear = "clear0";
defparam ram_block1a0.port_b_data_out_clock = "clock0";
defparam ram_block1a0.port_b_data_width = 1;
defparam ram_block1a0.port_b_first_address = 0;
defparam ram_block1a0.port_b_first_bit_number = 0;
defparam ram_block1a0.port_b_last_address = 2;
defparam ram_block1a0.port_b_logical_ram_depth = 3;
defparam ram_block1a0.port_b_logical_ram_width = 8;
defparam ram_block1a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a0.port_b_read_enable_clock = "clock0";
defparam ram_block1a0.port_b_write_enable_clock = "clock0";
defparam ram_block1a0.ram_block_type = "auto";
defparam ram_block1a0.mem_init0 = 4'h1;

cycloneiv_ram_block ram_block1a1(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a1_PORTADATAOUT_bus),
	.portbdataout(ram_block1a1_PORTBDATAOUT_bus));
defparam ram_block1a1.clk0_core_clock_enable = "ena0";
defparam ram_block1a1.clk0_input_clock_enable = "ena0";
defparam ram_block1a1.clk0_output_clock_enable = "ena0";
defparam ram_block1a1.data_interleave_offset_in_bits = 1;
defparam ram_block1a1.data_interleave_width_in_bits = 1;
defparam ram_block1a1.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a1.init_file_layout = "port_a";
defparam ram_block1a1.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a1.operation_mode = "bidir_dual_port";
defparam ram_block1a1.port_a_address_clear = "none";
defparam ram_block1a1.port_a_address_width = 2;
defparam ram_block1a1.port_a_data_out_clear = "clear0";
defparam ram_block1a1.port_a_data_out_clock = "clock0";
defparam ram_block1a1.port_a_data_width = 1;
defparam ram_block1a1.port_a_first_address = 0;
defparam ram_block1a1.port_a_first_bit_number = 1;
defparam ram_block1a1.port_a_last_address = 2;
defparam ram_block1a1.port_a_logical_ram_depth = 3;
defparam ram_block1a1.port_a_logical_ram_width = 8;
defparam ram_block1a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_address_clear = "none";
defparam ram_block1a1.port_b_address_clock = "clock0";
defparam ram_block1a1.port_b_address_width = 2;
defparam ram_block1a1.port_b_data_in_clock = "clock0";
defparam ram_block1a1.port_b_data_out_clear = "clear0";
defparam ram_block1a1.port_b_data_out_clock = "clock0";
defparam ram_block1a1.port_b_data_width = 1;
defparam ram_block1a1.port_b_first_address = 0;
defparam ram_block1a1.port_b_first_bit_number = 1;
defparam ram_block1a1.port_b_last_address = 2;
defparam ram_block1a1.port_b_logical_ram_depth = 3;
defparam ram_block1a1.port_b_logical_ram_width = 8;
defparam ram_block1a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a1.port_b_read_enable_clock = "clock0";
defparam ram_block1a1.port_b_write_enable_clock = "clock0";
defparam ram_block1a1.ram_block_type = "auto";
defparam ram_block1a1.mem_init0 = 4'h3;

cycloneiv_ram_block ram_block1a2(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a2_PORTADATAOUT_bus),
	.portbdataout(ram_block1a2_PORTBDATAOUT_bus));
defparam ram_block1a2.clk0_core_clock_enable = "ena0";
defparam ram_block1a2.clk0_input_clock_enable = "ena0";
defparam ram_block1a2.clk0_output_clock_enable = "ena0";
defparam ram_block1a2.data_interleave_offset_in_bits = 1;
defparam ram_block1a2.data_interleave_width_in_bits = 1;
defparam ram_block1a2.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a2.init_file_layout = "port_a";
defparam ram_block1a2.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a2.operation_mode = "bidir_dual_port";
defparam ram_block1a2.port_a_address_clear = "none";
defparam ram_block1a2.port_a_address_width = 2;
defparam ram_block1a2.port_a_data_out_clear = "clear0";
defparam ram_block1a2.port_a_data_out_clock = "clock0";
defparam ram_block1a2.port_a_data_width = 1;
defparam ram_block1a2.port_a_first_address = 0;
defparam ram_block1a2.port_a_first_bit_number = 2;
defparam ram_block1a2.port_a_last_address = 2;
defparam ram_block1a2.port_a_logical_ram_depth = 3;
defparam ram_block1a2.port_a_logical_ram_width = 8;
defparam ram_block1a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_address_clear = "none";
defparam ram_block1a2.port_b_address_clock = "clock0";
defparam ram_block1a2.port_b_address_width = 2;
defparam ram_block1a2.port_b_data_in_clock = "clock0";
defparam ram_block1a2.port_b_data_out_clear = "clear0";
defparam ram_block1a2.port_b_data_out_clock = "clock0";
defparam ram_block1a2.port_b_data_width = 1;
defparam ram_block1a2.port_b_first_address = 0;
defparam ram_block1a2.port_b_first_bit_number = 2;
defparam ram_block1a2.port_b_last_address = 2;
defparam ram_block1a2.port_b_logical_ram_depth = 3;
defparam ram_block1a2.port_b_logical_ram_width = 8;
defparam ram_block1a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a2.port_b_read_enable_clock = "clock0";
defparam ram_block1a2.port_b_write_enable_clock = "clock0";
defparam ram_block1a2.ram_block_type = "auto";
defparam ram_block1a2.mem_init0 = 4'h1;

cycloneiv_ram_block ram_block1a3(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a3_PORTADATAOUT_bus),
	.portbdataout(ram_block1a3_PORTBDATAOUT_bus));
defparam ram_block1a3.clk0_core_clock_enable = "ena0";
defparam ram_block1a3.clk0_input_clock_enable = "ena0";
defparam ram_block1a3.clk0_output_clock_enable = "ena0";
defparam ram_block1a3.data_interleave_offset_in_bits = 1;
defparam ram_block1a3.data_interleave_width_in_bits = 1;
defparam ram_block1a3.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a3.init_file_layout = "port_a";
defparam ram_block1a3.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a3.operation_mode = "bidir_dual_port";
defparam ram_block1a3.port_a_address_clear = "none";
defparam ram_block1a3.port_a_address_width = 2;
defparam ram_block1a3.port_a_data_out_clear = "clear0";
defparam ram_block1a3.port_a_data_out_clock = "clock0";
defparam ram_block1a3.port_a_data_width = 1;
defparam ram_block1a3.port_a_first_address = 0;
defparam ram_block1a3.port_a_first_bit_number = 3;
defparam ram_block1a3.port_a_last_address = 2;
defparam ram_block1a3.port_a_logical_ram_depth = 3;
defparam ram_block1a3.port_a_logical_ram_width = 8;
defparam ram_block1a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_address_clear = "none";
defparam ram_block1a3.port_b_address_clock = "clock0";
defparam ram_block1a3.port_b_address_width = 2;
defparam ram_block1a3.port_b_data_in_clock = "clock0";
defparam ram_block1a3.port_b_data_out_clear = "clear0";
defparam ram_block1a3.port_b_data_out_clock = "clock0";
defparam ram_block1a3.port_b_data_width = 1;
defparam ram_block1a3.port_b_first_address = 0;
defparam ram_block1a3.port_b_first_bit_number = 3;
defparam ram_block1a3.port_b_last_address = 2;
defparam ram_block1a3.port_b_logical_ram_depth = 3;
defparam ram_block1a3.port_b_logical_ram_width = 8;
defparam ram_block1a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a3.port_b_read_enable_clock = "clock0";
defparam ram_block1a3.port_b_write_enable_clock = "clock0";
defparam ram_block1a3.ram_block_type = "auto";
defparam ram_block1a3.mem_init0 = 4'h3;

cycloneiv_ram_block ram_block1a4(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a4_PORTADATAOUT_bus),
	.portbdataout(ram_block1a4_PORTBDATAOUT_bus));
defparam ram_block1a4.clk0_core_clock_enable = "ena0";
defparam ram_block1a4.clk0_input_clock_enable = "ena0";
defparam ram_block1a4.clk0_output_clock_enable = "ena0";
defparam ram_block1a4.data_interleave_offset_in_bits = 1;
defparam ram_block1a4.data_interleave_width_in_bits = 1;
defparam ram_block1a4.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a4.init_file_layout = "port_a";
defparam ram_block1a4.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a4.operation_mode = "bidir_dual_port";
defparam ram_block1a4.port_a_address_clear = "none";
defparam ram_block1a4.port_a_address_width = 2;
defparam ram_block1a4.port_a_data_out_clear = "clear0";
defparam ram_block1a4.port_a_data_out_clock = "clock0";
defparam ram_block1a4.port_a_data_width = 1;
defparam ram_block1a4.port_a_first_address = 0;
defparam ram_block1a4.port_a_first_bit_number = 4;
defparam ram_block1a4.port_a_last_address = 2;
defparam ram_block1a4.port_a_logical_ram_depth = 3;
defparam ram_block1a4.port_a_logical_ram_width = 8;
defparam ram_block1a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_address_clear = "none";
defparam ram_block1a4.port_b_address_clock = "clock0";
defparam ram_block1a4.port_b_address_width = 2;
defparam ram_block1a4.port_b_data_in_clock = "clock0";
defparam ram_block1a4.port_b_data_out_clear = "clear0";
defparam ram_block1a4.port_b_data_out_clock = "clock0";
defparam ram_block1a4.port_b_data_width = 1;
defparam ram_block1a4.port_b_first_address = 0;
defparam ram_block1a4.port_b_first_bit_number = 4;
defparam ram_block1a4.port_b_last_address = 2;
defparam ram_block1a4.port_b_logical_ram_depth = 3;
defparam ram_block1a4.port_b_logical_ram_width = 8;
defparam ram_block1a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a4.port_b_read_enable_clock = "clock0";
defparam ram_block1a4.port_b_write_enable_clock = "clock0";
defparam ram_block1a4.ram_block_type = "auto";
defparam ram_block1a4.mem_init0 = 4'h3;

cycloneiv_ram_block ram_block1a5(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a5_PORTADATAOUT_bus),
	.portbdataout(ram_block1a5_PORTBDATAOUT_bus));
defparam ram_block1a5.clk0_core_clock_enable = "ena0";
defparam ram_block1a5.clk0_input_clock_enable = "ena0";
defparam ram_block1a5.clk0_output_clock_enable = "ena0";
defparam ram_block1a5.data_interleave_offset_in_bits = 1;
defparam ram_block1a5.data_interleave_width_in_bits = 1;
defparam ram_block1a5.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a5.init_file_layout = "port_a";
defparam ram_block1a5.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a5.operation_mode = "bidir_dual_port";
defparam ram_block1a5.port_a_address_clear = "none";
defparam ram_block1a5.port_a_address_width = 2;
defparam ram_block1a5.port_a_data_out_clear = "clear0";
defparam ram_block1a5.port_a_data_out_clock = "clock0";
defparam ram_block1a5.port_a_data_width = 1;
defparam ram_block1a5.port_a_first_address = 0;
defparam ram_block1a5.port_a_first_bit_number = 5;
defparam ram_block1a5.port_a_last_address = 2;
defparam ram_block1a5.port_a_logical_ram_depth = 3;
defparam ram_block1a5.port_a_logical_ram_width = 8;
defparam ram_block1a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_address_clear = "none";
defparam ram_block1a5.port_b_address_clock = "clock0";
defparam ram_block1a5.port_b_address_width = 2;
defparam ram_block1a5.port_b_data_in_clock = "clock0";
defparam ram_block1a5.port_b_data_out_clear = "clear0";
defparam ram_block1a5.port_b_data_out_clock = "clock0";
defparam ram_block1a5.port_b_data_width = 1;
defparam ram_block1a5.port_b_first_address = 0;
defparam ram_block1a5.port_b_first_bit_number = 5;
defparam ram_block1a5.port_b_last_address = 2;
defparam ram_block1a5.port_b_logical_ram_depth = 3;
defparam ram_block1a5.port_b_logical_ram_width = 8;
defparam ram_block1a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a5.port_b_read_enable_clock = "clock0";
defparam ram_block1a5.port_b_write_enable_clock = "clock0";
defparam ram_block1a5.ram_block_type = "auto";
defparam ram_block1a5.mem_init0 = 4'h1;

cycloneiv_ram_block ram_block1a6(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a6_PORTADATAOUT_bus),
	.portbdataout(ram_block1a6_PORTBDATAOUT_bus));
defparam ram_block1a6.clk0_core_clock_enable = "ena0";
defparam ram_block1a6.clk0_input_clock_enable = "ena0";
defparam ram_block1a6.clk0_output_clock_enable = "ena0";
defparam ram_block1a6.data_interleave_offset_in_bits = 1;
defparam ram_block1a6.data_interleave_width_in_bits = 1;
defparam ram_block1a6.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a6.init_file_layout = "port_a";
defparam ram_block1a6.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a6.operation_mode = "bidir_dual_port";
defparam ram_block1a6.port_a_address_clear = "none";
defparam ram_block1a6.port_a_address_width = 2;
defparam ram_block1a6.port_a_data_out_clear = "clear0";
defparam ram_block1a6.port_a_data_out_clock = "clock0";
defparam ram_block1a6.port_a_data_width = 1;
defparam ram_block1a6.port_a_first_address = 0;
defparam ram_block1a6.port_a_first_bit_number = 6;
defparam ram_block1a6.port_a_last_address = 2;
defparam ram_block1a6.port_a_logical_ram_depth = 3;
defparam ram_block1a6.port_a_logical_ram_width = 8;
defparam ram_block1a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_address_clear = "none";
defparam ram_block1a6.port_b_address_clock = "clock0";
defparam ram_block1a6.port_b_address_width = 2;
defparam ram_block1a6.port_b_data_in_clock = "clock0";
defparam ram_block1a6.port_b_data_out_clear = "clear0";
defparam ram_block1a6.port_b_data_out_clock = "clock0";
defparam ram_block1a6.port_b_data_width = 1;
defparam ram_block1a6.port_b_first_address = 0;
defparam ram_block1a6.port_b_first_bit_number = 6;
defparam ram_block1a6.port_b_last_address = 2;
defparam ram_block1a6.port_b_logical_ram_depth = 3;
defparam ram_block1a6.port_b_logical_ram_width = 8;
defparam ram_block1a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a6.port_b_read_enable_clock = "clock0";
defparam ram_block1a6.port_b_write_enable_clock = "clock0";
defparam ram_block1a6.ram_block_type = "auto";
defparam ram_block1a6.mem_init0 = 4'h3;

cycloneiv_ram_block ram_block1a7(
	.portawe(gnd),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(gnd),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(gnd),
	.ena0(clocken0),
	.ena1(vcc),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(!aclr0),
	.clr1(gnd),
	.portadatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,
gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portaaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,data_a[0]}),
	.portbaddr({gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,address_b[1],address_a[0]}),
	.portbbyteenamasks(1'b1),
	.portadataout(ram_block1a7_PORTADATAOUT_bus),
	.portbdataout(ram_block1a7_PORTBDATAOUT_bus));
defparam ram_block1a7.clk0_core_clock_enable = "ena0";
defparam ram_block1a7.clk0_input_clock_enable = "ena0";
defparam ram_block1a7.clk0_output_clock_enable = "ena0";
defparam ram_block1a7.data_interleave_offset_in_bits = 1;
defparam ram_block1a7.data_interleave_width_in_bits = 1;
defparam ram_block1a7.init_file = "ifft_8p_fft_ii_0_opt_twr1.hex";
defparam ram_block1a7.init_file_layout = "port_a";
defparam ram_block1a7.logical_ram_name = "ifft_8p_fft_ii_0:fft_ii_0|auk_dspip_r22sdf_top:auk_dspip_r22sdf_top_inst|auk_dspip_r22sdf_core:r22sdf_core_inst|auk_dspip_r22sdf_twrom:\\gen_natural_order_core:gen_stages:1:gen_twiddles:stg_twidrom2|altera_fft_dual_port_rom:\\gen_optimized_memory_delayed:dual_port_rom_component|altsyncram:\\old_ram_gen:old_ram_component|altsyncram_obt3:auto_generated|ALTSYNCRAM";
defparam ram_block1a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block1a7.operation_mode = "bidir_dual_port";
defparam ram_block1a7.port_a_address_clear = "none";
defparam ram_block1a7.port_a_address_width = 2;
defparam ram_block1a7.port_a_data_out_clear = "clear0";
defparam ram_block1a7.port_a_data_out_clock = "clock0";
defparam ram_block1a7.port_a_data_width = 1;
defparam ram_block1a7.port_a_first_address = 0;
defparam ram_block1a7.port_a_first_bit_number = 7;
defparam ram_block1a7.port_a_last_address = 2;
defparam ram_block1a7.port_a_logical_ram_depth = 3;
defparam ram_block1a7.port_a_logical_ram_width = 8;
defparam ram_block1a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_address_clear = "none";
defparam ram_block1a7.port_b_address_clock = "clock0";
defparam ram_block1a7.port_b_address_width = 2;
defparam ram_block1a7.port_b_data_in_clock = "clock0";
defparam ram_block1a7.port_b_data_out_clear = "clear0";
defparam ram_block1a7.port_b_data_out_clock = "clock0";
defparam ram_block1a7.port_b_data_width = 1;
defparam ram_block1a7.port_b_first_address = 0;
defparam ram_block1a7.port_b_first_bit_number = 7;
defparam ram_block1a7.port_b_last_address = 2;
defparam ram_block1a7.port_b_logical_ram_depth = 3;
defparam ram_block1a7.port_b_logical_ram_width = 8;
defparam ram_block1a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block1a7.port_b_read_enable_clock = "clock0";
defparam ram_block1a7.port_b_write_enable_clock = "clock0";
defparam ram_block1a7.ram_block_type = "auto";
defparam ram_block1a7.mem_init0 = 4'h0;

endmodule
