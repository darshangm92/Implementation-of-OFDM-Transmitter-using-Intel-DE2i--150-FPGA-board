��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����軽���S8��A�>-?�������p��a�sx*|���~O�JC��'��l��Yὥhx�(���������	͠�i�+_C��w�pУFVf@v�r�Q)>�4A��B�x��lcU�w�ƈV1��!r����>h8M�7/��8o�ɢx��K"��7��\��x�WӴ���b~.=ave��$Z�rG3A����ш[�ԕ���_�%�0�t����y���D�eO�%Ը���Z��?��:6P)hRJ�;��E��]�b��\��2[�U�K��7H4��Vb��Z��no����Q*�栲�|_	��S�WO�g��JF?O�:�����:��5�F%F��v�k,--�w&����;�aV��$ ��z�3�|D��1bH�4Gb�O�.�~��(�uwZw��� �%�����}v�kW���H
<QĚ_������hG�!(dWȜg�^_�����!��f��p]{j ��g_��P�w �FB�z�c���빧�Hq]hRO��2�c1^$s�O��z^R8���^� ���z^��I���()�ٸZ�Wm�+��=ǅ9(d�t���?� "�XE"//��ΨߥH�_�6Ѳ�墓�
lJΆ�֟�ҏ��������[X�(Zo'b�m�W���e��(��q�.��g��#�N���A�w��*ů����	7|?�<c� 	�,�\]��e;9M��4�M�z�e�Y�.DZ�ۚ�o��9D�p��)Ɔ����fP����Qi���oW`|u2#�0����s�Nq��Z���͐m��7UB�Kޤ��LA�1�S�j�/'�q���'�����p�_Z���y�Kx��}�!�<���e�IFIW9�qM%
���x�{`S�D�,HJ��H]�L�g&�!Vi�e���f��TLZ��Hk�6糀�Rt7oc̡3�gN��>�*�K!oH�(�
L<�J�%Ȣl�{�-��(��t>Qw���~AڲA�2$��R��q��������� ��%T0T�4�l�-�)�O�b!�w������m��A��Q�)Ovz
F�U�꯫�081������z%�7Y�Pu��!҆�R$C�1'�\n��T�~&�r'�x��w�>�C����=��\�:Gv%u�PF�qQhyj�כ{�
�#�)���w�ن�+1`u锥���e� W�)�{��*�7 �p�����7�.6�	-O���)�i0�{�}"|���T�7&R�F����K��u�
n=�+���	|f���@O
X�R���(��`���-���'��d�[�����tw�5����|:�i���~�+*�8J�0�_�)�K��0��	W���Ѿ�d1B<I�JU�_��&�Q�dy���q���0#.�Q����k��N�vI1�`W�SP�kP�U<mn��;"	�B����p��S}%���m�l�#r_~��܌K������b$%KKW�Lt��y� Z]��Џ]y	Z����ѫ����ln��PO��-��O��n�7��2�$�6����Ȯ��I�9�W�2�i���7ɓ����0�y�R�!U�u~������|��`#���Y���o�go�"H�N���k�fCpx�4���'�c<[�Νl��!ob�MzYI��(�˘�e����:-�&0�9�F'�,' K�D�+����}̦�+�>����-�8&%S�-�����:�{���]2@Y��/�wm�u�Z����x���I)��?|
t�X�A,�W��8�k�!��@,��V�V�5=�6����H�C%��-^��|�>��)���v5�߆��}Hƕ�/���z��5
a�={�g��{�GL�Z�D�{%i1������x|Ck'u(k�dKϱ�&j��^.4q�\C��U�v<a\SR�|o�~�����c�8��0)��9!ֱ:|�Hڐ�7M������@"��A}�e=��]S������Aτ]ҫBʂ�/\�WB�4�����"��Nn��|���������M�j2��.�� =Pq�˫��+�@uf�k6��!;�-�U�Z!|�}h�C'�����S;�9
A�F�́���{6�<�X�췇|z�&��s�]2]�?�Nm�}i�*��7���c �����`]���x�U�ki[�CA�k��(f�F���Rg�5np���X�!f�W͟
R�Ԙ�4���ŋ6�hQ׏�?d�|�|��=`e�=��.��}~s���{��/=F�\�z�;Tg͆
�>����		�Y�X3ĥ��t(�Yd�����#���~���o<��O��"2����3tu��<�E�:���MJC���^�U�]p�;���+���\��_2#x���5�
�i��C�׫�##ۚ� �Nز��}�q;�&/�]s>���$�q���z$S��U?qԶu��h�ë�ʳ��b���C���=�jcIg`�k;�q��2{3��XB8�zq�71�DA��|n�� �W㕢�W�	t�;N�4���\�B�(������x
�b8K��r�E���L��̢qnb�N���sȧ���6����7�R,(ګճ�1K<��Z�}�����V*߻hl �7����\���;WK��冪���TWsi�<'��'ż�W޳��aG�j�&kS��h,h2ʑC;Ƶ"# ���o/&�|yJ/\Q��w+�Ťq�޸�Ἂ%NzH�O��w��j�L0ى��-W��٣I63m�B5�9yn��.t򇐬��QP��G֬�h<D��@���Ǿ��HKQG�z�*��I�jF�d%B�^ѥ��hW�G1(�]2�����	G�1���I�xK�/���B�����f+����r�*Zwݺ_Y��+�
�� O��i׾EiQ|O�pb�'9�Q����=����H���a��
�R��İ��]�X��;�v_���ӹ�1>������Q��wJ�X%���[b���Թ�T\����O��< ��?�7*�,�0�|D�VBt����|��Ͽ��q�@���4rGU�L��e�SB��M�b�n���6�H�2;7ƀ[��#	����)��.���1�h���"dD<�ȳ.ݤ�Fl�2M�qչ���%Mu5@ �߃��܀�-�|4�q�6v��ʒ�+��|��4bjy1��§�s~��ͻ��b��R�l��m�e�3��c�,�.Ա��M_i��,����d�_��\�ݼ_X�d|B�\��jn�非�e�SLK�\w�ɓ���J�C�m����?�ꉶ�Z�����K��=�\��B{�k�@����Z.�k[@c�^^{xk\9'X�9�L��ڞ���:E{J�R8����9��/CV���f��8UE��/�{��z>}^w==���������/sԁ�Qn��WIi6ډ��V���fX!�DQ���x��N���w��oZ7~���T?��Os�h5�-O"X�@X����7}!����.Ԇ�!����e^?���Sc�M����>�U��`;QR�o��~z�
��`���Uؖ<�U"�gw�{@g�LL16��/��T��q,���|r��Ww��\v�������:pz�?�R@��,6��#�D�����9��_K�ԍ���K��PQ��y�u>���Ef'6�5)DT�b�}�|���J��Ve��v��B(����/�y�`*�,kĂ;/�_�Mv^*�Ǹ��C?��ya�;�p�
b,�����5�d�s�l��yDL�p�~�g_�MqlV���N-^NٽRGyoTy� ����"G�~1Q���l�����9� m���cu�.�l�Ը���ܠ������ms���=�#*���%9��A�r��]=>�_�.��Mt���PT��f^V;�����(�$�؅���h��b)���>������(ьB��^Ĺ�I��,���9�Bj���S��g�[���"dطs�<j�W�[/�DN
�����kVs�`T@�v[o\�j�]N�e��Ob��#��kT20Е���H�E�>��BNH({I!<F�Y�g���dr*��#T��3�6��[^@�laK֮".OVy��Ք��]sxft{ YJ�Pl1Y���!�Bb<��%N�9}��Tr�I_L�ޔL딳�lP�M+�:)U��
��ESv�-�VsQ�T��\eȞ�/~r�0����,}?s�[]7������d?��o~�M�l�������(��m4���*�Z��iPd��(�>b�b��=7c�,i`�.�P@ąkr�K)#Tn���	�x�V��[׶}��0��ͦb��9���pj5��lE7�a�`;]P�z�w�y��y<q��n/���������Z{wM/�Q@�O�8�mPKG�� E�$�и���?�j=ײnL7����¶0���*܉ ��=�#O4mٍ4�c�j�L�b���q\� �*~�o:�}�ʳǚֿro3{��s7�x�=Wd6/�5%��`��+��m��T��t��y��Cp�,��b�s���sD��o ���F3�y�x�
Iy�m��0	��������W#t�A�	C�+��gf���f��,�j{d��e�V��0��N1,)���s�@��ZZcכvf["4}do�_�ج���tH�O�8g�v�FC���)�;��$"��ޤ�3���p�$N���xet����!��j����a�)���n�Y����,������P��(/����x	8�A�0 =��l�'��8TÆ��іr�F`�p�A������O3�Q�M�DdT-�W�x[���m,>k.(�����4�ET��n��
�&�[!��.
�Ix������&`|���O+��v~4*��gQ0ڣ/d�����Q�T���a,���q:w�fH��3`�d���'�%�����U�@�,�`,����n�<)��kh?�(J%g�/v	oCpT������Hl��PE#1���!�#݇�7�])l���B��K,@��G�?b!�n���z�3�����r=���ERȥ�a�/<8�eP{��n�A��fg���S��I�Dǜ��?�Ҳ�Y;D���H()"�
���	8I��S���Q���%��H�}��l~nl���׈l��s�vM��U�#'?���*�_?��)_�I�9��;�<�i�$"H&�gY��K�x��}ѷ&�U�qK483M9��%�����M@yP>�*��Cn.�;�ar�NAvzC���j�h�"�7<t[K3�U',�݋�W� mUOF��{�z�91s^_#E��e����0��K�ߚLwT� ���të���~�����cS��LBAȠs�����Q��&i�葁��~Ȉ�7���b�Nկ+�+(ҹw�Ҽ��M�
?ꘪE�'pO� V��RJU��<���2��������r��3�i�"]���,�`�J��$fNί����x �w�g�c$��jUw�p����}_���~'�D�o*�c��(|�&���o츛�K����=e��F�M��j�N�$n�J�&������aV?�f����f�(�r텑]��S�&k�ީ��X���>�4�x����I�$���lbd+��k�B�b��5���vkO0$�ɇ��� JT��s9��݊E
��W�>��ۭ%+�W����Q)���t=�B�[�f�%�-(3�N�rh[�������:( ����&�P���׆(%���vE�d<�$��˞���%��-%����Qb����P�@�����D� XQi
���R����yJ��?���?�=h�gj���wD���9s�����U_?HU�; �'g�Ѿo��#T�<�,h�HX���J؝�p:^G����K�������e�B�(K�.kj�&i�j����ψA<�݋5UGàP&}m�Mb*�&'��Z�~�O����x��D	 �07��V+�����	�x�
������t�1Gf��_\������Ue���ow'ۗ)O��xq�Q�u ��0���򜻝p���EEąh�q�D9�X��?M�R����2L��p^P���$0�N�)u3Pq�U���2�ke��$Y ����U*�����r>b�U�3 ���R��V��D�)I�����k�ѐ����&���i|/��:`V�+�R8�E<f��v�����~}�� �~���v�ѵ��7En
�w߇2Wv{��9�U�\o���@�M����Έq!~�|��@�Lh(,}-�T����H��RE��M�;� [oq�KWǮM��/� �y�}�؝��(�ݬϕVq�>���x�G����[����>�B��'Q���A�i�j&󙧇�Y�[����
il�D)%���~�
:���P�T!�kD��,� ��ұ�0��1�HK�͑����|�ज़�m�*G�U�p}���+
������Y�j�y�W<93�7���T�%v�i���i��NP@ϰg� 7qYW�.�O9YVc��$is^���l���1>>�!ɘO?G=!bp�̢Pq=i2(����g�rC� q,��<�#u�i)����[Ȟ�M��Ǣ���B��,J�<��$[+�L֛e�N�{����p�b_����K�(㗶������>���ʲ�Iꐝ�>�xV��R){5��	(5�O��Aȯ� �qA��:�'��������uL���L��<�e�������TfII��=P2�<Kzp�w�>��f��	eߦ���RZ@^mx�Jv=/᛬DW�1����Bp<��O���[Б�O��C.���2� z %�$�RY�׶�GjP�d �{��nDe�	�S�e�O6���2B��(�F��X�h����h���vI�&�#��e�ÞP�N��%��:YAG�a!��B���\g�e�/�X��J��I�?�n('VB����rs,�e�c� �6�+����O�C�ھ\��K��[Z^;�
	%������,eSZ�.+Y�����]^�Vu=�q���q�jQOf�}Q�����[a�Zi�ގ���28��j�Rpg�tda�����ɟMX�"������˵�X#l����{�������;Y�{ʈi�;����$�y��Y"h:�y�Z��0����H\O(бE�%G��\4����E=�70H�\��j��%r�=�	ј`gf�5����T����}�.^�=�˟��,���.2@s����v��h��4|���W�b��t��E]�ZKn�l�e�UP���ޮ��`���m�c��@�4#��>��BL�H�6�E,!��o��"��J ��X�cDl�H��+|q4?��Kى��	��<����J���t�7Aڒ@�^�r���r�3�Iu���>�p/5ݗ���"6�fݫ�c��Q/��T�қ���P�@A�D����]�S��k2)
�[�ȏ[Ņ�ho�Y3N�-�I���v+܃t��;�1��x`wq�(m�U���Y�qx�)�<�Ǉ.%O���ŵ�}ܝ��8eD��B�s�8��B�Qh̷Kk�E"/���ux/�`I�#�7�X�T|&��$5�>�>.����ޔ?�^��yIT�K�G�'����Z{���̑��m����*�)4@��)���l��>\
��*\U�ӊiqczzi��i��K�auA*�OY�6�T,ϟ���,�ʕYz��!Cfq~̊�pL�ؖ���{^�q���M��l$EypT�<���D�A���Z�G����}��i��NaT��:� b�}����3�a�Y�|������)�wHr�k��Vq*Y��"�ٯP��>zډ�+dy��������1�X�ts1��E6��rQ/�j�v�[jլb�v@�k�!TS��~�O/��Mêhl3�m&s�2�Jb�!�>��Π*�H&Bq0{W-pv�1�7�^7��ƒW]���'J���9fn�=A����d��u�7�t �y����t:q��`�B�Lj���*�b�$4kr�b*M�0/�\�-���3ڳ�ػc�;� 6��`����zq�r�����LK�z��m5AV�D�k-W�&x��K9i&]�l|d~��G�!0��I lNf4�˪�skC����z�\��~�Z��C�����_'�p���'��*��gl}�ң��k�ppU?-2p��+�UZF	M]*�s�y�jH��b#l�Q��L,F�s���[ֲ^���}'�7r��E�d6�Z���x�ȍµ�H�c���Ia�h;y񬙉Ȇ5�S��yF:ɘ%�cwTk/��|�|o��)����el�V�lج ����<Kc|{@|o�T�M�&�0`ׁP�\�L@�Z�*���B:��[¥z� ���AS��#K�KҘC�.g�]L�o�������4��W���:�=l� *\�ǲ.�G���vt�<�J�'=Sa[H�O���P�&Sm�j��.;b�����d��r�ҭ��o�w�[��xՅ�g�ݓ$���|��m9p����G�{,	��sR��&{��'S�띆W�+ݫo4�+Ц;㷏̀rT�BJ���%����}�d(�FZ��Zq�N���b�D���P�:a�a����K�ֶ�0�;L5,h��Is��ڮ�[ab�	Ly�(5�Z�d_�d�s{�j���cA�.����>2G6�2*����O�Wޯ��������0�2�:Z�5�p�{Mq�3Z]>��X&Q����p䪦���nָ`�.�S7��w-��vTp�ϻ
�sQ��BXWHI,C�M�
���V��.{���k�V4%���/T⸝�"f�&|���}�{)���}����;`kο3R��B�=S�gR� P[�^�F�ƹ(��MvD?ism�;����0W�j���G���Xy����3��m���^��2�H����rB$�[�<�;�O�ڒ,.��Q�kԼA���H�AUe��{^�xk�V�Iǝͷ����U��mU�6*�#��'��t Zt���ЁWy=2�R�����������9�|:���Ko��W�E/�Hu��|�p��{H�
~Zs�*�\���$
��_�qN�!`Y|��� &�0��Gd�H��F�?8�,%ԧ,?4u���{��1@�4��XL�Ѹ��٢Q���}������u���	����!�[��q�ZD\�r��(~���W��H��~x��mV`y�7`mdZFXJ�EЇ�� g���L�G'@t%��]���:�o-��E����+�X4�A@&sG�QN&������V���됊��ts��ף���V���q������\�lp�y�~l��yw2���f�����d2l����A���l�=�a�7<
��gp�@#lG�k�Q�eO����(#_�A�t9`�F8��zk�L&��0*�Q#+�R̅y�m�+yN��^�e�o3�4��KV���ng�\�#X	Iw=D�,�˄p��B&L��LJ�iiZ_-���ǌZ0��L�%w=iA��"	"d�D[�rJ�՟�о��d��N Jһ����mĳL/�hA��iqM��fR�V�\�q�z�y���$sp�V3���:�g�K�j1Z�l�G|��2��EN�v��}�"��"J�G� �c' nܶu�O���]�_�Q?�99��R����U�����|-�=�I��_ʊz�d$��OW*̅Y�@���ėwn�^��
�8�%/��t,
\@#�Mڵ�(В�Y�k(x[�=>���N!}k���C����^u/��I(n�ASK��s�V��oAw�4����|����~0"�~�,�\F�����+X�;_뻸�f
��~g өE�r��5H����-���u�j��4�ׄLf���Y�	��Ȝ���;J���.$�ˠ�d��{�Ʉ?�,�A�Dͱ��R��k�:��/ѵ� �oz�7z;���^�7F���4��n'.�E����@B��"���t[�j2�����b�a�����Bl=w��G6���z�W�����YL����z�pHwEx蘞q������ �n�^���s?�g�����U��5��-ZK��J�-�ӓ�Y������p�hNDK�|B���Gj�2���g���:y��m��ۄf��" 'д�h�~���m�~��6mP`�'|Ȱ[@�`Euͭ<-7
;����-{��Q-#��UaKDe/�#�/��+��o�A����*7ܯ	r~���K�Z��_I��J[�=��]h`���)��L�BJ���u6��#x�k��v�W|�[�f�a���o˄ ��B4��Mq���(�>u7y�S��d�J��+!m�Xb r����<�1/QSU�]>)5J> r�1�c^��I'qPpA�����p��a��
�q�2=��^��|)˟�q��:uy�1��������5��1�n����?��Tl�&�W�
����}5�� u���Df�F��!���+�V�7�3O�{ %���vl���G��{DG�mq��1c�|�flW��~ T*��}몑��G��/I�<�~�r�ȍ}z!ms�cA�Uɿ�j.���L�;�
�~+q~�����^*�5趐Bj5�4��v�c�?L,U{�1�24!QY��e�z�'Z�,��֕t,�F���T28	O&��s��
Z�o[Ƶ�*���y��{~�^�˚,��W�(�j�O����jѠ�_���H�B�vU���=��pƟ�-E�F"ȍ!��'	��H*ʴ5(� ��y��q,�b�t�)����h��q�m��7O���4�#H�B��P��'I�q7���o)�%ם��(ԩm'����&��a���d�8�����N���8�i���Ѭ��H�<:�h���V9J�@4�e�Z��8}���������lZK�$Fu�b�򔡼
֞+�}�����@0��Y��7�کa��"� E��O�0Q۝����Ƀ�\�5��Oӽ#��nBd���'�5���g�d����8��ڔ�{�"&��K�KR6����i�:@��F���L�#�Zu�����!��?!�\40qrX�6'oN솕��Z�V#����^G&#�(�H�z�D�,���]��Sͯ×�=��g룱�O˪g;�ׄ�Тse�3���1���:P�a/+��D#���Dգ��܀5�ʕ��o�J��ԐYk��{ �z!l���z3-���(dQ��x��l�1���V�҆�%(�N�}ע�y�/K��_0�'��!�T�m0ηA��QM����/#��,`{��]����rs�r��]� x���K�#t�j������j�-œ�FD�̣��wUӧwa��Qd%�)ȸ��S�n��鬝�8��Fd �4�ϻYB�x�\�7�g�����C�W�(��(Ƃ6@(�$nC�uՀI���n�ԃ���H�Pj�"�mI�s����{�<{5��ND�,m�4�n	��I�e7~��9m�Lr�1�K���Z��Y���Z-5s�����B����$��t����s�:�=s4"� �_�^�W���F�1�@���6~��B�Ё\�a\�<%2Ћ��gNG򺙓����I�R0��j�cJ+�9�v
��BZ����]Ev�S�҄�,{�
BD�jp}DV�ĻJ��z�ȥ���ߋ:�	яO�w�>Oϱ@Ѕ/qy�����k�Ϫ׺��Q���·-�o7g�Ap`�7װ	�o��ɺT�;��Ep`�_���ai4��ްR�w���6�EL�a��O��P�2����|�u��$�d�f��O�/x=�O�9`���c� �ʏ�"/<�.�k"��sP�w�r���N����a����ܷ��O�[	�2a=�F��a�
"ì�.2H���g���ޙ�{���\�6�v�B�,�I��%�B�&�v"-���hA��W��NK28�-#��IA	���?�H�w%��?kA�`/�i���sn��di����F^�Z`��Ĕ�!�d��9J��%�V&!���d>�ry�';ޖ�5��E�o,�m�l�#q���Y.v��~G���"�����/� ��Sy�4jB������h]�R)��:>x~�|�_�7�
!���^}��j��,�.W��]���#?�1QU�w<��$�U%ȶ��P����:�xl�/d�粎�:��R|t��V]��:w����K�|����f��1�Mm|�Ä���� q �{F���R)}N����㥞^�Z����L>����<I� +F���rcN�7�N»�2�6�$���w�	����©��dkB�{҇D���:�v	J)]~�:�:窫�֓�@RkZ�$��x���0�T�{^]�\v*]�h��v�J_-X�Q�qi�nlo^Ҝ�#�� ���$�����^�B:*��V'J^�,P������%�NS�\ğ�\��rU��#O�Z�ЍK��?��\O�j�i��-d���+A=)2�؀F-4~D�Z�����#����Nu��ԉ�V���.HY�+u��Jn���z�� $�li`x���G*�p/ۂѽ�@�&����}!��c����z0uk"q~1Sr/-�#�H����?o�<���J���qRx�ڶx��@*��J���� ~�'�8 ]ykh�Dq��@��d��Ө��e�:sW;���,��g�&�T�.��(斑�Ey��йXѹ,��(�|������~�p<;Pv�&��bk�Q�n���:��]��%��Y��B����&�0��k<Q�Z^�?�]`2�&_��o��Ngq��$�l�<�:lJf��zZ�+p:���Ǳ���{}X��8���#5�% h�'���qb�K~#K��ʠ��i���5s��� �J��mRG����{��ǁ�$^܏�D&`^]�)|#yMAɠ�gK�Ϧ�D�(�����'.d�}�U^����Z�U�C��8SCބ���yl�e�D�
f���x���s@R?���{kd~l

#h�,���`���;��Ʃ
7fd=��[ z���gj-�ufTF�]�1�5��}�j2���&Vp�`v��J�/�4zZ��S�6w�d�İ�B�Y=r�O>R$��;�M����.�+���!�&�=�=y���Ds��`#�i��}Kͅ���)R��f�|�T+��Uek!����&��P4g���C����>�eX���i�c(���.kO�J��O�d'�,��d�՚^��o����J�m�>[ >4�O�2�^���j�ĺg9�6dcn�����f���_�.�S��5c,<�(�O:ޒ����UAU�X��<�yc5���@���)T���R��ɮ�{�)�Zc��CE:���T��U5D��UP���R���ѧu"82��2�Z�����2��|�B_86]�c��Y�K(!N�~U���4�ER��Wy+�Y�>���Ņ3�y-VЗ�Q��'�E
Ha��MmZ���X�`=�xr���f7��e��09(E��b��P��7�0M���x��A�Y��s���+�*w�r!A�����a��)~�ǲx��`�P#i��iZ~�̤��n��`gFx!UC��M�k7���&��&�]?+��ߟL/	�U}�O�TGf�Q�ƶ;��2eŝ�2���;u�O�41��u�s�
7dKY��/ׯ*��H.��鎳�>�nMn�\��jN_�g�ٌ�ԳP��0�v�.�Aq֞Y��&������	�ڋ:�E�_x��]���44!���΋�	�(��b,����/e����f-����#uT�,16te�`��h\R*�{�p��?�9�YB�!�����>L̴D�"�����S0d��6�����W�6O4�����1���g���M��<j%�줗�s~S6J&]��:|�`�cH%b�#��w��`㾖}r�^�b�3����߲A�aUe�A$G�+[H%��h�k�d$�4��#��wC��"��,�J6�1µ='�e���5��\x�B�I�e���mI��6U�n����M(�o�T�/��j�o�B>�����9l��Jg�ػOAWJ��x]V�V���b�@^xe�^�B��N�0�S������4=�~w���/���oK>}jJ���JGG\>���ܴ#Y��/t�����Z��;��*�'i�5��h���D#����`���P���pu�!*�J���_��%��7LE�Yr������_��-b~i0�:Y���5���z��8H�V�Xg U��c~�I�=���T����a�>�6
EyטVԖ���l�F���㰭�~�i��m�I��"P��D�Z1{&�]����Ћ��5l��(?�lߧ�����-C\�@>�+%F� C�t���@�a�H�@~���礥v�F�q�'��%���V�J$�	�:.��.v�Z- �N���I�h������*��9��4�����hR?�,������M��o�+#�VP܈�dcu�!��_tH��i�/5*�p>�ó���&�����*؂ahi�w! `tм�����d�M6���ҽ���4�� j�Y���zD�p�n�I`	��f��I�� R�����{S�:�jY_��ѱ�)8E�x�g��.��.tN��ږ��"��=xY�O����%���V�����K�G���-E�~{߀!>���9T���ǝ:1<��u�De89�&��3����;���BvY~a�$�r6�=�ؿ���2�:uJ־����WΌ+{�i��Ґ�R��/\S�Lh}O7��ᖡ� ܹG�2�N]Xe9��a���u�qC�Ș�A- TP�Ƹ�ԑ��^}���;��	ўn���L�u1������P����4���'d��ӊG=�|��1��I��QO�>=y4e�n�*]���T��1��^RܵuX��z��d��'��HwP5��2��R5�������54jv&g�J�d�����*K\T��|�Oݑ�C����RbO�!�D���+j���#cx��"�O!���Px}D���i%N��*.�3�+ۖ�i%q_5���.�P�>1K��Q���P�Ű����T��[ڪ��� _���$I(��$V;����B��}�Cx�T�+�m���n�T�+9��+�JV�J3NJEP���r{'9Pd��q�8�׌�Z/8E�`�*Ɏ�Y�"���餷��\t��{w�(Ú帆;�v�_�N�'N�F}��0�����Z�J�!�m]�t��M�ΰ��]|~m,��!ۉs����<n�l!����j?�kY���x�����vPKxU����	悤�hT��a�G_�+;�K�:j�#�.�Ik܆49|��'�����^-d��R��c�*� �|�3�30�yOq ��%e�*?��ϫYx��J�T��٪0����ɶ�Q�;���℠��Sr9���91l=r"	1 CA���He�|^Q#`���x����>~u٭x�������/��3�u�F�4G�I����pc�|��>�D��?�М��-�?=U�}���`���-E��jNZv�צ�D����9v+�3�?%�s��E��@���Q�ʋH�����	���E��Fk���l��+O��A��3����Ƭn]]]��&�Z���'��¨�bv�o�[�۷�O�Q�yR�l����Xr��.�˛1���ۣ���~˶�iq�������`Q7�zAw�ѹ6&}����[p��������0����8�VT*�aM�r�~T����Pi{c�=D�	�Q�1��C�&�����Wp�?G�lQK:���N!xL	�;�|�ŀ�5����1��(3��e���GlE�wYB��Ng^��e�����+�#�ʠb}�mE���:�����#��c !�F����{'p��@����#6Jh��?&�1�FҌ~甽��u�d�� õO�)9���G�u��D�|������/}��d�oD)rL3/fJ��"��gm�����nSuv����l�k�ط��32l��z����-�yĘ���锆O�eS���A��v��
�|��N*S���:�swH\
���ܡ�˛�8��K+�}�`�������,��x��	j���]�B/�C౉�.���U���XOm�P�{�ߕ���{�Y!�5#�*6�P�$�6����"Q��`4'U�w���.���˰�$u�te�uW�S����dި�P�R����?:;`�6n
_����l ��P���G�����J��E�}7� xM�'.�NGI��y&}���'����N�)�����՘zK�X�)���U���L!%���i�������)�� ��Y�Qۧ��iZ>�f�0�#V��\x��1HCgA`�� �a0L3�`���.hy*y1х�|8�
��lf�vu.�k�ę���� �&$� c_DI6�۞���A]�,�a���o� ��)EG0�a���n�p >*9rm��$�3<��ྑ�q�!�e5�/��*t>�.��{u$eY�`�<ԂA)?�QP�n+�(�9��0��}.�O��Q��^�&ѥle���R����r|�ى��D�V�26E[lhR�{��&�VT�
�0U�\���§�=�('QM��"��DU6R�vO�bB�9qA�'��,h&��o��d"��>ϣVgj����mvP�f^�1��`���I�h.�0y��m��׏z��/)�z?��9 ��t��jl���&�%�ݙ�;0���'�Ə_�Z}0��Xvԙ����,�9��1o8};��
S�"0���Պ�ު��]R��8L�Z	;e�o�G�Ԡ�Ѷ&�k�AY�" �`��d��l�Z�B C�?�h�]УRH�o�\�%�Ӻ�C0H���(7*	�O�i��ۙ�{�K�p��ww%��U^T�{����J�a6�M�}q�^��.ط���&|��d��B�5����:��y��QQUO�yI�@��H������i|�lyZ8y����9�K�ne�ʸC��r����Ĝ(��X���%`��L��i �nc���O�[|��M�';��	Q��l�g�ѿ�x�����<����B���"S�S�Y�s������E`&����^�0�'����@��!��TT&-�<�^�7���� 2kS(�N���*�S��w�xp��ؗ��?֊�̘�A��p����7�
<�H�1O1Hp$r'7v�o�(Byk��mM*fHM�-Qak�m(n����� ?�h�d�D�KV������\�vג�?$��j�J~V;4��pE6�:P��HF�@B<�-��ٲ��wƁZ|h,N�P��;���8� Zu�@�al�#x8�����+u���܆�k.���õY��{	SJ�Wj���^$���2�_0-"�,�����1���3��x�������?��x`�NE�q����	I#�8:��P��L�>�~���Ȯ1kpE �G��d-^���,��(	���216"�;�r��WW���d��^c̪��K��i�寖���\Ԫx���N��L�}��D�]�G�5 -�M����]�����W�w�!�xcX�l����f�)���ν1��JZ+�Un��U�K���Cl:Iӳ���.�Ƅ���=2P���>!�:��6\���P�v�k@�f��
z1�wD���!�[6�[�$qo}a
��2�1��ey�(�!���}j.�&��7���+���i�3ugjE�k�o���������%��j�b�{�z�S�Ҟò��FM
��^��Hg^�ձ�p/P���]І���0.�ͬC��`�9��|.�U*;���b�+�7����o�
Cb�-E�=�Жt�.�Y�yr��c����X�|���i��#w*tv��6MG��M�C��0��몤ZP�¿��R\�F������_[)t���&U�B�r� ��
u��a�H3���Ek���"-���_A_ߠ����/7C��\��kH�_P�9](eo5��s`I�^.��������@̍0���ź�|�-�b�]�`HĠ�?^Kp�OS �:x�����*�3���ͨ-���)x�#�k�g�y��~�8��ْ�tB�����Iq�v$������+W��b{&;<���Q�d��fg5J��IALS�n:}�@�k���E!''c��*eH��!��W��i���,�^o�]Ͼ&�hO[�s�25����S��]F��{�P������)�Isp,˗�ED��8��W��*�W�+g��`���ۋ�ݽ�/a̩W���oª�D�XWz�����c��Lo$���)�Y�ɋVlȝ�A�_Aw�]M/���xn7�e�i����ka�14)J���5bdk�h������k��9��^��/�A4�ZJ^��>.�<�[3;�zf����2�=����K=�߾�Ah)ի	C�%V��Z�}t�Y5��^��h�NndJ��p5j8��#9CP+�`�	Y��a�ܦ��F���[��r��d�������R��>�n��ԩG$�7�����ψ���TVh똆�g�5C�±�Tmt{2��y?�p��n�(�jzlr��լ�,7���.�[�%���䮩g�L��ayt8����%�ʜ�g/͝�]X�an{����̑Y��бi�J�n��q�	"���P�+��;�>5#-��qX�rP_t$oWa��$�A �����ک\��]|H�8���¼�=��}ӵp}-��q�6]Z�/�7±u�]n gM�Pv`�:m�V�b	jOF�뼓WOz�Ng��Br�_p��s�z�����(��q	]� @9��D��bI^m\$��9̣U�/��k$��l�|O�hG�[�~�o����t�����S���G}�t�O����_	cũ��:*�#Bf@�����:���+���GB��&&d�}bhM�<��� ��K1�)0�������G]f�mi��jv�v�,c��aV����L'����A��ق ��B�z�H �IC��C�'g��8(�u���+E%2��h��2yo�%Zw��=�c'b�+T��ִle�а��#�,s �M�?<']��xT'�\�'�R2�r��O�(�ÌC(%xt��t/*���/x|�3���툱�N@z��]m���	Z�]d�g���C��X��H>u6��t����q�D��a�Q��e��7��Za�e�-lS�P*����U�f؛��}z�����i$"���g�Yv�U�Ή��uor�}���j�#�`���m3) #��Qhm�;h�v~����;��VW���gv����{Z��ԉ���ka0
ɋ�cb?��Y�P�;q���v �S�8!���? ��#�k�ݘaY�%N~t�@�f�X���D{�I�G�6I����JX�g�;b(�\���;)��<L�j�}E���z�*>� �{�@��(�5�� �g3���~�Y�f���\��v���3P����KQ���7Yx�yv?�n��v G�d�I�=�l��%l�(	RT����u'���엽t�L#~���WN��p�3���Z���#�8����
��2�C�8U�T�F*X'K��T���n�ɻ̂Y���vـP�:�$�1����{���8Cdx�p�R�ځy����"ꈚ�Z��d����/m7yw|���\��τny�����e:J�R�D�<h��E���0:��_��}6��5��pk��u:�y1�1��ٞ�;����/�{�bq@��$�zѽ� ���ӱ�؎��dm��l��a��?T��:�S���ۨ|�D:��e��k�	����ԣ5���Aj�8���̷���m�&p�D�.�Ѵ�������0J1�&���#��xD��dE�[��6/�T�y�K�!��K_yb��!Z�T��Y�^e��7���ջ�9Y�5E�X}2,Q��+;Ç�&�*d+0X���y�]�@��(��$[9�잱�T��R�o�K��)O��5� ���b Tyi�ktL�eq�v���gk�	_8�/Uej��͆Y-�
���<d�Z���5�d��M둈'e| c�N9������)p\8��ϻ��:*�C;�!�F�Թ�:�D]��v��H��zn��CǊ�uP�b���	���'Y��	�Ɗ㷠�;N�"�zHOh�4.��\���k���4��~���%�'l�H.�{#u��)��nw��ݙL�tŬ��]�-�^Md�:�x.��b�ܒ7{#)I;E��pi6n�x�%�UKh��)�o��p	�O����L4~�ac?��P���Zɛ(���E��8/4�ON��j�F�v�ϼf"��󏕄�
��G wuL�P��;07Np��8��4ԋr1r�s,R��	���0p58�*8�Z; '*ZU>q^ǎÿ<�ׄ�6���52��+��tӖ�u�Tv� IG�B�Kh�ݗ��=@#,h�d���γ�	��}X(�ĂF
~�@�y�9��]� J�o��)o�鄟�/����o?��vv����a#WX˴�n>0����I����3p�ѠB�p4�m�Π��o>K]��U���@P_r��X��I��Cf�����h�z�M��P��R�H�����v�r��*�	A̓Eqe~�*���{]��bMI��b�l�H�R�4�6R$��f��!�Ρ��I[_S��k�_4����T��&�ɢĜ)2�f�o��S�����}g�iJ9�vZ@{�,$�S�P]Tb���"�swV��A���:m�lN��=�l�X�}�Q�sK��kvO�H-�����/�!n�EӁ�б�N8K�J�����v~4�sYO��-j�-9(WLK�S=��u/` z����j�Z]���}�-��g9����_H�=�
�mȗ�����:^�D�-b���S�=�6�ҿ�`���*�cn1w���q�r�.g�����b��"�_RLP�A��-4��ٹ��t�#|T�+C����GTpZ�0���p�S?{
�9��p�ۀ�/HN0���7�=0��'��Jh��v�� �E�r�ͷx�� �Z!����#9;E�{CG^�Pj��IxWW�T��1�Ȯ0E6q��A�4��g��Ͱ�v����ꈻc�4�]@�e�螏���'��/i�Վ�G�M�>�}�6��AK+m��GNE� �W��S�9������'���၄s��r��Aq{��۹Fv��M�s��!���{���Y�o��4����e��?�Ϥ�H8q�3�]t>X����-OXL�!�Q�cًqN<�y�+��Y�F-Z�e] Z��-+'��� j�R�5��4u������|�9h�����"x�����ҳ��I��O���Nv�����,���ռ(�Q����J�XР��7�c��qX��	!��@��gQ4��a��\��a�<�~彻���>��;�7c�x�ڌ�Go�P�ZK��Ҫ~�~� ��,֯��#)/�Y�(j�� ��<�<c̈́�o��/�ЃK�����+4�ٱ�fïա���.�t�XCQ�w�2��pzJ��smf��/��0��I&���P�G�5� ���9�e���+�/�z�\�y߁b쬇><��3x��M�;u���r��<&>q��J�B�X�	 ]�kM�:��|{i�Y�C/��pZ�0~Rx�+�fR��A�j��wi~�_�K�@J�)����O�8���[E�O�O�Ep��C��X6\�`w��p׵��$���f���d�D!-��uyE$�R\�W<��M��_/8R�$6��"��A[�,,X�H�|u�� Q�
��%�JiB4��x��,��e$Wh���@q�t�+A�}9�ޓs��3�È�,�x�U(����NN�z�ޟ��6(���0�0M���>M���M�c���m(DP^�ߡ�{J���OnkQ��P�s��Щ6�	�%�K��O5Ю�F��ܗrF�G���/~Q7�UF��(�S���=(�o����:���=\��Ce��xK�g��l�b dr�����m)[9Y�4�!�\����Z�p}�5��Db:+i��T��Ag4tq�n�@��Fݲ32Km�*Q}ג��~��lˁ՟��b�(��#��E]I�8�dd������n�e�
��x�oB�2���X,�SK(��8v٫CshWr��e���ٳ���������ɢ_&�G����Hpș��l)��C�L
S^kx㢣N�Q�V2h4cZ4����2T������ɣ �<�ɖ'�/��<;(��L8�����uL(N�s��wbj��`��)kj�{��Hw��	�&�A������f��p�>3�{Ӛ{D��fے�.%Τ3���b�&,���g�BE)���+�a��d)!;@��`���x�Q�m�H�*��]���{��������t�a����;�%�*`�U]����T�@�`]4��Ap ���ް���sF�h8C����i�+m��u��4�f�?b�O'S�[��0L�V���h���#�IS�>�h�$������{A����k�U�Ӵ�-���=�@��Wޫ�RZ��0o����������/1��Z���b��R�ؖK�:��m�y��#r���Y�C����!o[��En&.�#�$���������=�;����՛�;��Sb��) 
�)�v��J��0��~<;��\*�A3�}l�ġ}틁�/��]	���Z�y�=_�J8v�Բ0��u�	�?��7����r���u�luoU���<����%S���h�w�� I?���`���K�O�2��U�P�Ux�(Y����#]1���_��~��p��Z��ï�3P_A��K%1㨖��c5jߢ`_�~�uttbf���t�\�Wى�̀�1R�HE������N\�L���6�K�l��qs��!_��JYX7i�"��1C����l�)��6
�n��l^�s��<�En�{%D��o�����ۿ�����Uxl*�@�C0f%��SB�}���v�Yꯞ��Q��#'6�X��I�P%CV��F˷�ɰ����
OT���}��`����7�#���_z�����;�M�\bR&G���/D���l����+'5�	�e�k�!�Vd������L`8~���;���@"ܓ�Ŕ���D��d6����0��.�U�v�z�~k))���M�9��]�
U:���ti��pGg����q��Z�;�8C7m��	i�a�G��G��;8LJ��~2�A|\���n��	 ��V�Q����3������ �@��#��47%B|�G�j�}x�����E�6���t�S ��H",ɼ_o�ϰ�=f�����Uދn-O��T�j���Y�?O�TX��i���ԁ�d�R��6R|������@��GS]�	����?Z2���y�b�b����.���GỊw^♒A{eΫK���я���z}��N�h�ᒵƺ'��M���Ԇ����S'm���P�a.o�3�%�!1h훀F�#���Q�~¡��H;=*�Nݚ�Z>G9�<���N�JN��A���%F;-e��ׯ@+�6C��rb�	Ck�b-�y���U��fX�H%�
�MՀ�f���9�b��ۊ���v�m4ǯy!k��VH���s.�o=���da��`�w1K�vA�Io��?AQ��F���'�Ac��U�<�ϧ
�����W,��E�`�_Psɡ�d�
��͏3�����2t�V��v�Z�/���:�ɾQ�yF��.�#��m���]���4{|×d��v�m�I�����Y��md�+]h�,�ظi�Oƀ.j_��)����T��:����`��o�,������5ה_��4��.�m����<?j[N�+�.Σ���!֕B�u��m���u��FD&HС f{��l�%�EQ�z�D2��{�k6Z��O)���E���&�Bl/-��R�6��L�`�mA��mW��lc�Y&��©gl�̞�_�[��Y���^�Αl����GU���ueJFY��H0�[SRC����a�{\uT��^�����{�A��g��d%w�x�Gۇ�\��-n�y��ȍ�[��u��*�U� �;��o�N�E��j�x�8�1�=�ÿ�آ�2�ɑ6̮U�;kR�I�e��g���L���SA�,݅d�%�/�pL,���y'��$�E�FAR��{�][�qA���=`t�ה�pӸ\${�y��d��:4y"M���N��uv�e���ð`E�x�8��G�BΟ����t���FyC���Y�V��u�:�|�������2i,����W�4��Ƒ\����&f�i9P,#�5�Ch��^j?���:� �}�ؔZ�B@�F�K3ΕV�FV-e�g�rKq ��X`B�fܽڽ��P��}������nN�$V�����[ڥd�ƪ�KO�V�Jr~u�!#���_�a��HL���#,e.ٯ��'V{A��k_@��\&U�|mr��Zp�D���$C�XEp���¦ځ��1���A�Q��w���$R6�Lޞ'4�9�$� [�l%�mE�� ��⊏-��3���$��Юk�2�+���N������`�!	������Ր�,�N�rSF��ƥ�fL�z���̋�B�_��3�՟;L�ą�/��7a��.�����Cn��#O�X�O�4߇������̇��]�ڝ D0	G�-�,�[��<�k�_G�.i�"
9���4�e�5J����/a���"U���J_w�s[�������q|.f\�\�/^O<Ußg�Ym�FJJ�Ũ?A��E�-T3fCZ􂚮�u�5�|��魵D���·�(A\ѽ�}�&�-����,x��ݣ(7�Z�#`A5�\B}� Ђ�׉���G�I�
��s��;&���Y�����$�h��tP(CjU�ܢ( Ð��v*`QpS�����݁Y*V��#\6QyY���s:Q@����Ժ'��K|5Cn�����N��ݧ����ڢT�!�?ǥvQ�kB��FO� �7g�������5��A%\�&W�v�=tl�P[����oQ���Z��ܷ�KG�`���[�h����橂v�
�J6������Ћ���\�s�u�@;��MY�:bzėu�6�ԥ�
BD8\�b�G!�Hg�/�߶����4׳7\�n�I�w����f��M��u�L6���Hѭ��-�W�;����^���䳶[Gp�R�)OֳL8j�\7�%X�h�nh��'D@�h�4�h�|yb]B�o6F\�~m[[�ip��,��oUB�,�:C�k}�$�H�Kl�Y��"���@`�N7R�	u��o�zM:d8 ����?Oz�Q��k.i�[��Pw�s/@����L��7��/��g&S�u, 3�LbTD�T:��,�h��Q��E��X�P�?0�\�'R�w2� ���2X�ٴ̭��'��Y�"��S���yZo��zů�Nm�K,1� a��1hn���(�v��<m3QtbDT�B��%A3�!��(��@S��?W�3�B^���,@ɱ���%�(r�z�]B�v��8ūT�X>�`�?<��Y��3R0� �M_gO�i��Pm��D��� x+y<�7��[� �W�����)�Ա^�h_	LWNű�`���є�pk�qzõ�3p5��r���������h�3WPR���s�����I1I�u!��u���~�����I�,����oUD@I��nիu�9K����u�Fp�bq3��B\I][�@r`�,���>����g��#���p��Qܕ�5�өDC�h�F H��/ɶ,��b����VÑ-jS�*O�ki�2�ȴ94yو�;��k���γr��qQ�uF=��]`M�F�GMl~2���T�U��+A��0�+8M��=�a'}W>�?׭Rߥ��qр�X��o�T(���s��Y*��H=x��vf|�
�����X'2B�1��D_����>�I��U?�#�s�>!vC.I+���G*�_�d�� U�o�U����|;/��uژ��+Һ�X倠�І�ø�e�.���x����5�8ŋ�)N�Ӷ�ƪ�~�����C��y�$��2N�E0�">s\�A������JE mV�#�Ζ>���)r9���6B	T9֖�-�*���}��a�*�<�~F8d��073�z���M�0��+*�� �?y�@�M�j�6c41���NI�g�J!�,[T��iŎ�!�Q��L�H�\���sQJ	5p��
�4ڽ~�3�QB�l\����O`�-���d@xy���,=`�"K>�n�����s� FM�`�I[�����Sr������.�WE�XC8�Q������������&AoY=Lߏ�%OpX���M�~����d��U��NA� �gx��_��I��Ye;p���;C�C낭�|׏���I�s2�yw��w��Q�:�w�u�YD)Rm-S�fX������+R# ��3�?B=O�͞��Ҋ�4�$�X�:�aa;oq�[1������U�H9���g��.��ևi�4e��qq�^*E)�f>��~_�	+�~��C�{�I�hU�9�DdPE�[�t~�_h�K�^82�>�gA8�����tA�����҆>��I�X�q��иQ���tx��F��iVvr5�)�Ȟ���,���W+R�<�h4??Jk9��q��3r
���Я)/I-�-�9Y`��l1��_� s�86���`�n�y�*�0�l������%x6E7�-j�=Eڸ���o�+����Cz�5��ٛ
�.�(�VJ73�ދ��ȞQ;�j��)|`� �M,hⲡڐ�~4֒��eN�t���pu:�N L��΢`F$��k�AV6z2��t�
B�'Fc�
���F��r���м��\���@�qEjc�����޵
<C����dH�Q����Қ��u���ư�3��c�oT�=6r��:�u{U�<,�Q�f�1k{��n���e�/G@֋�OY�}4G�-3�k���t��"�]<��X�����T��W�s�_qꨌ����3�[@(n�<J$
@T���	yJ�%������4�[��P�0>�Ck ��,����u}�zWp���ȑ�p��NZpsF{G���w���2W���ơ���v'�(���S�/���<#kvaZn�����ώ(�x�BY �R:������M\���w?�8TK��K�1�#C�r��^<��0�0�>��ߥ4n��;Vz�L�-���]}��@�BԘJ�7�v)+/�$��]���x3Djdxh��إ�N^%o@D�V)b�1�MK�}B	�q@2IX�PVmX��׾�C*7�BѸ��C��]y"� ��3�Nv�i�B�?��>�d�y��{��Ԃ<S�Ɇ�yF�Uz�J�0�JJ�81�5�m�D$��l�v��^9f��l�|����!+k�g�MnBXw��
��7�)����L$��#:��4`��% a��bƏ���R�&Li����6GMutTM���c�eD�O$��i�j+/�j�1	8Mm0C Azh���ijY�i��u���{ۜ���%��2����]��f3�͔��X��"�Dc��%-fK۹̼�a i�V27�1{'%�8��NY�4R֥Q��9(�T�����ٓB�5��A=���7�#�C��.��UuDrï�.��yeyV��r���(Y������R�cMV�n8�z��c��s�A�گ�4^�-��q�'�ck�f��lﯪ[OKl�^=�]����z�o�|zx�}$�c�
���P��
�)�#�S�� �o�2���F+Y-x��	?���'裊�vE#ECjjh�\,�K�
�F��S��o�N�В1�%�wJI����I���|��l*w� �m�E�5z#G�a���Y�'�?[g�Vݾ�E��'���vC�y�N���3x沺I��F�<gIY������mTY٩��K����fC]��!`Z�c���U_W�s��'��x�P};S~i��E�a�]��|�Ę��f��A��BT��Ţ��1�u�D���Q<��5m�?���F���L
,dY|���;����� 0M���3[TI`�?ֿ^�9Eo$��[�'ܬv۟���	l���`Ҁi��.2�VK��oS��
�
|��	�jwOcʇ��-�K���bӢ>۹�}Я4�FC\	��i$m���VBᙅB89.r� ;�����j-�-ڐ�swl��m��*ah0ra�:{�D���\�����,$m���KL�b�_��+U���vE��puL���rwҁ�Ì#=�'C^3�������sM�1?�75M����#8�QT�P�Kx�����ʖ������EZFշD^|���;���c�o��431f�0�R,��@�-��z���+
m �
�J�r�1�L��~��h Ykߙh��<ɕ���u�Nʉ
Y�u�S���|�}��B��Iyٝ׋_��4�/,�ɂ2qW{�O6�V:94Ŝx���.SƝybB�:��F�����e�1�/«=����Ŏl�+��M[T��O�2��L��V���tp}s��U-��6
q-z�h:=�)����Ϙ�9/��M��Vʇ��߯�6�c[����-�` �A6�ٛ�j �Y����g�߿}IZ	P.�
�>�*lq)�������Q�(]ЏCI	3*�50��k\4���s�"�s�#U���@�#��H}x}�!����pY�_�}�]}�,_$~U�&���O�����9���)m?�*�T=��ʗ��^ ����얪2bf�!Q�j� <CA%�1'�p�� c��f$��=3��/��h���r��w�����\��:�IU�� mZ��%��*l��U`����[�/��F�D���Q���XF��uᯘ�t����d\�v԰��%����ra���[������p�p� ��4��PT�V���66Y���[�-��u�5��vA�CK�Ag��f��ʺ��aE�ns�m39 ��x�5�9���G �����a�G�L�D�=�� ݴ���?ԋcV+m~pla���d:��p&����¿&�$����N��4�Tk��9!Yt�O�bgK��{#�Hƃ)eEœ:�amm�`�I�������42�	L�+�H�����I]�$d����r��^vd�e��GJ$��:�M�o-��T g+u_j����N!�����:��S?S�'�L�_qR�x
M�b�g�%>M���"��
�M�)�w�F#�\\Ouf���~?�᪦��j��-! p�/�����'�ݭ��o��)-��XXy���p�w��m3 �Sy�$�����<���}o��nnB%Қ��&�������ש)�_G�����a��xg�M�;���B�t�T#*��Xq�D���-���ZUI�3�Qi�V?5���Y��������h�*`�ܭ�(чy����R>m���r��{�lBvR�s�>���,��}��v]��,�a�/���n����{� WQSq�сO� n�$<�ll-�g��&ʨ���2����ӌ՝�V�w\�~%)r��tG���+2��S���μ��w֕H�N)��r>S.�m�7}]�p�5<%p,��A��-@�/+࣐�"��`�B  ��􀆻�K��7�J��g��TA2����g��["�UR��U6֜%��|��' ���g���qB��B��NN��g1�#�EH�cP�RX?�릟��Sb�h>�M�*��x.�:���U�/m���!�I^��A[��y��4�2�a��p#���Ei���S�Qj��f�Y����m���W�Dݡ��F&���&!fT�[����� ��
ݮ_���̽0h���2�*Y��B!���&H�c2A�T��Eˁz,�p�
&E�bl}��ɽ��o)���Y�����mz~�G�C�i�����#�0^�nS��#_�׫v�i���1�h%��/�Bk��AG��(a*���;7Gn�!j�#�<�}�ڏ�X�G�kn��I�*�)~K���Ld?�&�`� E�y_P�pg�ܠ�t�|������'��`�+�31���~v�+�ؖ���| �ǌ�d�W�Gg>�\��L���:��T��9.:�^���H�Mz��mj�<�+�uehg�*�����R�,2/e��GX�7���!PG\�)�)�$����Av[�H�������]���Y�<.�����%3�:�uE�M�8A@��۩�8,W�N�_k����$�8N�>5���Uv=9K-�b$B�憙 \�����$�����^T��[�Ԇ��6�C��H�c�i������=�
#�B�["��g#�Q�������¤�92̘I9������k,g	:�Ԕq�Q�
�
Lx�`ۀ�����^�"�����n��P�&���T�X�V�3U��&�9��S���e�NGC����$���d7�����|�ohg�Ψ����m�i���H=V�K-ܪl�R�_��Y�<T��g���&?�r`ń�R���>��:��r�*�QݣM� �=dDp��R��u�(�G����7����Wc��f��>�Է��0����6)��&>��~��m�F>��2�z)wݥ��ɨn���YX~u\����r��P�?��[�*��6���P]K�e�v��eFz!w��`Ζ�w�l�CT�0���7%��YՍ'@Z����ud�vV4��,��^��r���	i<�W��mq�a1�}���|��+7�q�/��n����@Z��z-�t���Z������ ���!�����l#����G�bD�䏜�{��,���/�!On���8 _�M��,4vA��� &@;݀��S�fy"=4��`IeC�n�L��
lV�؁R�g�U��'�˃W�[v���_9m� _i��:��`�±��:/�5��c��y�t踐$X���?��GO�������S(f����7>�"��,1r"�,XΛ-�1�Z��b}FB��!=��6Qf@w7���̨�Nű�t�\�&^�qc��[���{cegyY���CQ#��N��F��	��o�ZȬ��H�o��p��K���ڏ��ڔ��r���3*�)�0��Y7���~�T�7`��������m��U1����f��w�_��[�-�7��:����{dU�A�Er�J!eE� ���K7%�ȫf���;7?��ۼB�ե�9�/�ԨC�H�[}m�͑``y�F�aF�2�%�q����D��Kא���o%�-K-�t���u�mK��[��pJ����R��Q[�
�����4O�I��=wqF����֢����S
�*��C�@g	?�2N���\UUB�w��kK�J�R�ԡ������ �{����E.Q�I���e�kt�/_r��ɞ�j�ܤ��k�.�o�5u].��:��W� J��7 ����;G�B%Iϩ���fu�����j�'b���.��w��q���/ZlR|p�JOӮr8[�`���o`�������@��OO(�j�K�Upυ�R^Jl����#�^�Dc�.�(��ܸ^�7��f�|��g_��rKZ�nu}�u\_��k(L������������fl��BY��gl-
����`kBг멋��[X�/�e��2AX�Iv3h���q�1R�`��uO�g�pm�6.zc8�����xG����k��MF
� ��|w�(�#���������)g�L}ۦ����d8�xp`0C4m�4�<8��ԏ�'TD���6^��D�y��b�F��X�ff�I��"�39��|�l�7�hq���9�7{YPܡU�+���X�
*K-]6Xo1�i�g�k���T��-��;
���CU��?��$
8xV�{��}�~�@+V3~���<X�&�g�'[G�x3�Q�s�͊���n������ ��I�/fp��[��Kb�2�����<Uf��_F�6���d��ܑL(�����f{��������"���R��ˠ��/z,��ކ�]H�(\�۴�6L	�EH!֞CثP�S7~���ɡ���������XR�@g�s����(Spwë�rl�	�ݞ�w+־h]�DD�=b��K4^q.9�Oqʒ6'dr��������%�ɧ�QAEO�i��=�a���F*�Z�ls�@��Z�V� �h%���(XK��S��<�4ֵ��˷ p!��ۭ��d���lui`.	�IJ�Q��]����>DGM�9J��o�7:�|t����g _�Z��\��a�¶�C٠�RXb�}Ŷ�LTS����Z]�H+�U`eF8��BHX0�@�.ja����Q��f�u��,�O���U�k�L�ل�:LYsR3ӉU�"y(]u/7�$T�T�F$��ёsɵ��
Q�i3h��<��n�ql+�g_=xee�F�`�*h<ˏ�OԸ�i��m��L�p#l�ʳ��8!";W��5#T.~S��`��!
��S;�S��d�\�fKaJMl�U�[@)����W�	���̑��wfB�M���H�zDVځ��ڨ��4��"?���QU?��H��e0
���Q��.<��J����Փ��5s0c�&ߤ��Z�xx�c߳Fs�K�Ҥp�
"���B3)q/��~��j��ѡ�X� 	��&����IUuO�m]�!��I=z)�@��53�T�>>�����?��AN�����/پ~0;��h���F�v�Z:L��Qu�<�������/n�ҙW&T&~kdha"˶{CɯP���tC@�>��^�C6�����v9<DG��'�H�`�m�����/(p�`Q������΀uH�s|C��m2,��e�Ք�U�X�
�����^� �nM���f]�	hCW��E�������26t��B��59:�����iB��/�dq�NTw�����e��w)~o\�dU?ÏU�kʪ���븕s�_�َ��rm7�I�)��
��0f
�5y�p4ۃ�s��ףF���V�G�R�,�M�M[�{A�G�4��ε���Ė��k��\.홝8��H�,�hij��yy�k=� �"��/Jl3i�ĀيG0�i �����"]h��3�3�rv5v�o݆�	J��sh�K�C5�][{����d���*�ᥦuP�K�Ö0���B����8�P�O��72=�ʻ��e>���s\:l��o�{��6m4�|~��V��8_�m
jcMgl}�6���N�w]z�X��Z#�:Q��ҎԪJ@q����f�rh������%�m�J��8�˭��S��q"ߎp����~݅;Z���iT^���?����-L�1��3�*?��!���9�p�F��=���������Boõ�uA�\�r����K�ؼZ셆6��=%�E�Q�Nj�:W��t�H(/�އ��b_�;����$W�=|�d1��X���*��mC�{_�t�-���&�|Eq�e���]Ď�Ѯ��>/��O��!��r���5V����nw��q�編(��eL���ap�A�g6?;���-rH�T#��0���@Yrd���*�L*�=�4/��Ь8�-� d(9��඙�`��~�$L���,e�t��C$}�`�QA�)BհWGC�Z���sk4���'2ֱ���{�{���nL��<�i��{����o L*�!D��m�&����120�t���v��/IZ�;?�����~NS���PT43��).���2|�`�=>��aZ'��P�ʔIn�� ��4�;rR�#��צ���Q��B�;����Ν�E���U|p�0�R���B�qV�+����	�2ۙq�w�Uw�R�F�|wI�	���o1k��b���F��5�v�s��,�t�����F�t����9�ͩN�Xf��q��At��ǵ�L���}�t��/Z[�rY2�j�@t����#U�{�M�~��p��ot>���,�BV��t[N!;���#O�S=��HZ���ެ�-������5k;�-'�m�����/T����M����؃8�Vi�e2��0�,-h������"�����!�H����xr��a3���"���;�Ӥ=<ό�W<J�r����� v�[)�V{�b?��ߚ8�
�M�)+#�#<&��ͬ�h	��_y,IЦ/�D/�	n�Cu�ۥ�r!��2+�9YcL��J�FXa���K�^ұ�\g��;Pd��w�[��bB��[�)�u��u�]���T�La�ʳD6K�<qG2��C��~k��D:�����_�x>Q{�G!o��c�ys�ZЫe���yG1��u�0�SάJ�ϋ��~Е�� ���K���*�~�t(�Q=���ߏ��Y71�����w̿!B
i�p�@��"7
S�K%�Q�@[��V�	$#����ڂv5zo��(]�j�,�%֡PV�0k���ܯ�w����$��_�5��K�-��þt� sE�=��>%��=)�g����|j��K4A �Y>e��\b�ր�q�Sߨ���)�kf��3?�T�=O(,��"���e�� nS�3��3�용�>���ٕK��t�FZ�����j�>��i"]{B����1��.��\��	LSc��,�7��C�,J���w��A�;�?n�ng�]�τ$7�;�!k}T+N�g�h�$,#�CC�1MQ�/H��U�������d��F�edʐs�e�����q��7ِ�����Z l̐g���ݥy����b�J��7C����P���<<����W�D=��!�ߜ)<4r!K}�S�9�L�?�\�2�`�ꓽ���M�Z)m-P+<k�_'���f�y��ê���ea	���tqi��fS��.���v�a��t	Y�Sp9R5aY�9*cH���t�=Y��D�=�ML�X���s����(��Ȩ���������!�fۋ���!�����_M;NOe�".��F
{�]U#�e��A�V�#'Á�2) ]QkCYb(��1l�9��`�����w�F�$�[��f���i�� JS�eT�`R\1����qa�<S�+9?�8wC�y
r�ff�qI��$�-������)�#ꮈ�:T����js>җ��v���X�?�}����:�[���5y��yQ�1u� d�tn`�axpe�樲����B�d"�o��v)�{kp�kw��3�v���u �ߋ���WXmŸ��7&�m�`���
*��A=_�Ki&����lM�#��(_��r�4b=�1P\�t��t��=�b_m~Q\PoA�U�*���@ ��|�?���Uk����w!�'|ҕ�φ�9q9霻���(n�4`uN_��^�����9�'��(�I�R*���+%���F\��BE����82G
Ϫܛ�)���>��`Vp�+%�ɱ�W�A���-�ގ3;�-����r��`\�4�KP�����DU�� �k�P6�{�(0�Zl�� şT�<OcR�S�	�ۺ�S���Ci�3�+"=�q���@jǆ��%��?QE�-� a�a@\�����.g��u��q7E�;��.��na��ְ������R�Q��X��<!�o�^F*Do��P�����Έk!�x$N�����'�l����'^�@�mDc��FPB]�m��!1heT���>�u���awڇ)َ�Re�A�&��O�^Z���mߑ1���@�Q/���+U�~��-�Qf�0/\Bz���>��1y�6�Qi� @�fFnV�/4ɟ�(}�B.la��}�x�����&L��]?8���0��^�D3uz��l�r��m^�`�����P�G�c�9��/��,#�;���q��$)x?�����'��JEl������!����}�X>oh��t���m�8���P�DAWP9[l�C�30ɦ\}(���Q��;;��� ':�X[$�9vWSZ�c})���h> ����;�����T^����t2���#y�T㽿�K���$�v����F
?u�`�f�d���զ|r�Lt�w��~���8���j۝$^�BE� �"�a�U�]jn���`�������Ƌ��;ѻ�$ߋ���QJ��H)��7ͣ�~u ?|�8� QJ��,u����`Qл(����1��E�=��ˤ+@(�l� ӥ9P� X�l��,i��^������\ W�����k¥ck2����u��OH��U�*�8�x��x�'Zj1���� ��'Չ�i��	�dg���zæԝ�`MZ�
�8�0i��w�e����Dǖ�=�
(?��"��^�/���)�rn�z���Uǰ�Q��KVu5�y_��4����ju�qqV�2:��rb��U��E���9�?*�S4��4��յ�L�H�"S�-l��Á�.�r��n��������B{TNOS!���El�\�����
֌�"��*�=��$��"M�&w���/��� ㉖���	A/,X�ic�$��R�.�������ba藸Kza����k'�Q=��0'�a��Np�fO�V��G1��H�_�p_�vJ�҉xC��!��\�Jh�jN����nW�`�J�d��������F��f`Q���ͺ��vD`z7�+I����RY~R�����Yܴ�E�C��øy� �q��[?�fl�l�5�
�=��6��������mʡ۫�7��s�#�tk����W���]0��2%�R`%.&Yp6�H�1r��,�j��"�%��
�^�A;���*�	�!��F�6�4~���x6�c�_�B���>-T�����X��BΥZ�H�c����hG�z�|�i�o�1, �+����Ch�=_�'�ƘlXTg�������"�I(A��*(;��}/����)�&�3 �Jh��KM#�~����j��şS��ɳR.���\ő=W97u�']}�Ml{.q��[�[�&]����d��D�c�6�诳���b/,�R�MZ/;�-�����c27����=��3s��Ρ#�Yvg0���Oq��Mf���P��S�@�b j[^k�ٹ�-k�Un2�#�ĉ3�;�n}JϤ>4�1>d����7Iex��r\
A�P>}!�݅�Z�� �Ȯh׹��ŋ�6c�g
Ө+Ʌ�W\��0ʿQ_3����#�\nE�Ep��HE�硴{)ҧ?+	"ř�M�����i���N�k/�x����͏N-��f4v���g�2���6x�SDp�?|k�At�@̌�� ��_g��P�J�E����<B�����Q-���J��!�X�&�/��ߺ�1vKL0��+�y��i�D�c�8�}��s�^���^Q������&VH�9�����Ӝ��R�
��J��b�P�{�l�ܛE�ǔ�w�n@���\rC�M�{Jl�T���D�����cEf;?����<N Qg�BLH��z;pL)�<��x�+�����r�����
F�'?s� 1�	 &~����8��~�f��_���w2�16�nyhǥ�$�[nC���eKdq�LF%�A���"���$�X�?�L�����l�<���>��u/�|>M�F��$�N�1��a�q�K,��g�x�ܜ\��(�*��a����V����s0kD��M�YL�'-�ن���걢׻C���|6��R��qx�n�0����K/t��;����$�?է�ʷ�}(�«��{�m��,XM�`���'���y-�gcRBNi�믩�j�X��҇�R��1ߍ�(,�������Iv~�Rl駘��d��S��	�D["�e@{#���Z��;�������Z����&�钪�E���3@�+)g�dm���0<		�/M�1���.��w�-�Ш�6.u��1/�	l#�ז;���E�\{˚�h=�Uem%�r���K�zPgYlY'�Oj�Z��R-������3�z����g5H`w�L�f�jG��I�_�Oq�+�	�ґ��/�٭lűSe �v:ѡ�|R��[Nq��պ%�Ɛ"�tC�����RW`|���sCT �;���3�듟�>�
:�V'�S"#iq6��kP�~�p[�|ܣ"�M�z)��D o���M�퐜�;Dj͕�]]�|��Ӱ'���!��\bg�a0f,��,�2��sK���jd!����R��BBN����2irH����8>MI�p��{��!��Ɗ�����ޢqr���G�T:mAE�q,=;�s �������ܡ��Ǜm��z���::�vѧ�S�$q��U�W��:1䙼c-� D끲�fa#7]}>QA��h�hE+�L�欂�s��H=�5��t�]絛q�!��3��2�pkA�Xĕ�T,�D`7���,� ʻ��<=�39�<�$��e���~l�7�=]����β�f0�>q	�Ȗ2��z%K�+]�,_��q�lQN��U�'�n՘�etX��6 �[�#,���O��)��X�w���+���B���0ER&T��g���=��ܱ��|�78�^����Kӝd��c���R��M�*�A�8�*��l�����|,�Be{3֜T(�7$��n�xGΟ�0�z^��yS�:�#�bb�m��[����d�s���Ɇ�n-�Ow;@��3̴D��Ŏ~_N�vmlBe{c#{ҝ�ov�:#��E��!�"=���1pX��g�;�x��UW�5�OpG���3���*� ]m�8�zچ`)����X��`6q���ᳳI��,h�ǿ��9�T��1��j�P�ܒԄZLIv�W]��̮a� ��7#��8�zBS��D�fζ�G���4�r�8z�7�j7
#����=T���j6ܥ�[d"49�5��� �\Kv7	M�	I���;�; ���H+�@N�>������G�pу�M�9W�|���:yK2�'�J��ӛzK�xG��pv�H���SB�.�u�l�0NeZZe�^J'Z+O:��R���L�6bsn*����++���-$���/d^a4��rJ�o1t�2=Рx��^�fd��_7Oe�֯"��ۛztLK���|Ñ�k�l3 ��qE��-�!�7%��1!lt	�"A��֘SI��a��[�î�'�j�|�J�*�PD�։�kV��ǒ��F����lʧH�(8 �����x��Mc@f92=y\�n �!��@�	^���M��\e�|y4��P,�͝}���x�;l�2׏6��/��˙.���T�v��_�.���-}�C�YV,M���na��T���D�-�&�T��ɞe���N"�+{}�r�Bz<�Kc,�ze4��3 .�-�#�φao�<?gB�
��D^��{���"mJ�0
$E9yU
y�73���4�n��=��n������]���l�,#]�:��l�q�G7 &&�Qr��5��ا�b������wVv(��m�B|��F�
gf�p�y1�4^����VDK"��z��J`13�|8��m�����	r�	��0<�kJnog��b-�e���|��������w�2�R�zA{)v�R,�Xv(f���*��m�/�9�D�&n��`йq�D7���^�	�rH���q��ң��
Ԃ�FFFr�Z����O���m���P�R>ײ%�Ӆؚ��,���
[!f>��xR�䪙��h8eV@)k�Vݖk�/3b�:C�#>M��m�@��::���Z{�sXXL�qwF$�+;� �y#|���(�]��H��~f� ���s"B����0̔�tK�� �:�=�����L�,o"�͈l��������M�4��z9�U=�\�Q��PDCT�1Y	�y2*aBo3��������f*���ǩ���S[U���C�gkTcY���lq�pGWv?��Nb��;��	pw�6��#�����_�G�9���˲i��\��*p��9�5M��.Q7�#x����w����_�����d����YG�۵��+Z m��-z�ƻ��$�T�H����`����۰O~���ܲ	���y���!���.X��I��o�t�C�<8D�M�R�n�O��{��W�u������f��_V�F��@���p`5y�h�aPH��b��ye'��h��ߛ�ο���њ�l߲�g�[w��5�G�.�6[�^)F�Nr|?��Խ���ȝ�?���R:/�ؙs�eB�}�����h�B(���qp|ڇ���&�D�]�s{��&��,+{J�p�'WXҺ�,W>�2���R�A���k��K���ʹ�`�h]Q���.�a��sNf�X���:���co��-|�i!K{6��z��G߁ub\�71ɅF4���� �D�$�ߕ%����AJ�Y����QM9Jt�����������OY{�U:hb8mSt���ڛ�	�-V�U���5������n���nNh�rv��r��pT���X�b�e��KWFd��Y�����h!�O��f�?;<��\����v�)�l67`k���?�|�ݕkj���ف�#n��Z�#2GV�)܈������L/E�z���}���_l
��c���2GH������j����h��/����mքٷUa7p�0�hS�J�n���)��+�}�}H{fv��b�cb���q�hm�1奨Q��:8a�Ñ����ξ�v�h�Ҵ�h���V�h5�ĉ�ڲ�o��eZ`֦𗥭����*�H��3��#/E��9��i,��^����r�F��{��HCܬYgt�5V--w��lo����sB9.?�?���xs+���7e�
��C>H�W��������%hH[7� �Vb�t�w���
�<K��@�4}�nG�H9`T�m��ׄ�qRP����z�Wޝ�{ۘ�~!��_ ��+�-a]2ي=�#�¶��))j<n6�:������gJ]���%6�m�Q�^�IEnj���U�ܬ��m&���c�aS�6����U�X@�,�VI�3r� ���@�h	7�h�櫭��!��vCI��ҧ�mW��c���\�FTL�>zwT����e�'%�����qqX�UBVx5|r7��	�Z�ْ<����\�&�'�I]z1S#���2�#k��=�*	f�jؠr)X����{�}#�5�1����A�#Q�۞J�A����6(#=��I-�-˂��B9]�1�������e�%SfeC�+ ���e���|���^Rwr��)ڤ����Xp�&��L��e��������޺���Ϊ��������6��:�I���}FMV�]mc��� �g�����_���V�O�#�mRbE!5�0M��F����v()ڽҘY������Ս�Ȅ#��x�.j�\�����d���7?�Ͽf�c�N���C"��4��$��}�o3��\�S���&���u����p�W�
���ο��2�ES�f�B���.]��:K��kv�?���$��ar�3�@���,��5)�6��P��J��YQ0�|C�/!�P'mB�U��;Ѐ?lZ�,��њ�t�n=ڇT�"�C��d2����NG}U��҉��G��h�<O��K�=�1�V�@Ix|�q9�Q��}V�H&%:d�����;l�>e#���A�q,K��)�[���b@�`�y���� ��o5��*Q�K�H�4b)�#�v�����ԬLcF4�6�<2�"}�2�`E����E���"J3k�j�w.�ZG�]�[�͠zf�opu��,����d���%�p��%�y�ˢ�G���?� !���n�F۰ϢCW���]k�A�����ƛy4�i�o���46�Z�v �����7�ۓ�J��_��1g�U_uFU�n��3a>OB�����L��Ӱ��,�G�N��D�k1�H����n�R�*'�8�����Q����8Y;H�z0*�
�(�Cx�ߗ��R{uq+�j�'.S��t���L�����-��
�d��~�}c�]T��qa'�CK�7W�&Rr���5čɃ2\��zc��1���R�����;�������o�ˣM� �$k��=�.�ˆ�S�0��f�Ĝ ��wy�@��&�dD-�IO@�Py���`e�����PD��|�Tc�1�ĸiEs��c��N�~�Au�&�bxЏ�_�X�f�,�#h�4���D�]�� ��U�~�d�s��;t��AoAR�%q�Jj}-�Zb6︩�&	ߌ�����t��<5hP����A����P4W�G^!_���kL�/P�RM�-	�� c�+xB\(}\Ω# 㮵�RD1]MO����'N�� ��G�Q96�y�X�e��GB�HD�ǣdh0JR��t�a��\�����
�:�%�i���!����=M�K���h3�kw������7ٿ~�����/��E�&����Ř+W?8����6@$�M-[�2��H��Wt'�S�OIȪ?�Iz�aM@|��Ĺ��{�zcF����_xb�p&�\#�!H�O%����4�� :�j?��՘{���Z���;>�=��|N��	�UA�<��k8AO�8T
���y���ܼѮRRW;�������Ң�q�Xl��Ǻ�7;��`
%�Ϲ3�Q'�N0��:��;*��B�|�0�n,E���ԬGJZ+�u�m"6��BRe�r���1�� qv�������`�` ���#������5	��)����5\-i>��yܯr�����ɲ�-�˺ilj����WR�/��.+uQT�U��>���逰�bŭ��yD��w�$�s� [�������$��2^�cC� �WN?�8\@;��mJ�BM�5�V\�h�C:�+ �q�!�N�w@��p�Jn<���y�ԃO�;�ێ�Q�ʶ�^;���Г��Id��%��?�>��X�>�p��	�#}M
Z�53^�=��4c����>����Mn�P���ާ��
�Y����]Dx�k�K���l��3
�ǳ�s�UK�c,7Si~�$��ARii��@I
7�l�U�i�x�>�B�,
�����s0���h�o`����4]u1;��fx��������g�3bh�J(A����`�Z�J��y�@D��)S�M�J?���������k�_PO��5S�%��I`��CɊu������,�q�2���0�e�1�p�{������{��.�x��%)4��ж�:mX��G��S�ro��>���W�^��c^��J�ޔڊ��R�J��_���6K��)���t�kcfDe���鶇�����z_�G-xç$|*R_Y!�Y&~���
�*X��*lrT�nr���(��S��{$[3mV=�
�)Iߏ�ǰ9@���X���tt 	3jr�����b��j8�L�ac�����q�Yw[��hBVUf�-(���b�#�>���
�,4�J&~�$|y�&%��)˸�w�����`����P�{-�3K��m-߸x�O��gD����z�ܜ.�70O*�̿-6A�>����kV�i	�t�d�l��
���"E����Q�#ɩh#�J�⍙|j��q˶AU��*�E�2H�9�Q�+�X�L2;�qv�D\�`�U���,o4,7���1��}7V�����ca} }:{�0��AA�u{ ����k�SF�.N�'��x��*nL釘i��������n�"�;oO/�*WX��$5Oʯ�>Q��{�<�L�`JXcak!��m7�ɲ�p&�͛��q��ߖ�h�;K�g�GIN��eajع�ε�P�-���>lm��
�'��ʝ!��*�UF�Q��6�_�f��s�%���h��װ�X�	l��<�8,2!���@�`N�y΃7֭y뢼�(�Cԑ�yxE����Ђ��&���r�����o���/v�*�ZG�YDg;�Pz�/��I��\ܞ5w�o�)�4���Ճ��R���p������1אڨ���y�d�PLB?$o�H
z�{����2��W(����ӯ@ᅨR��}���	վlX�ҥC�UO�ɡ���0���,tB�	�p�O�����J��hc���J%�i���N�_gK꓀�%r���/ܔc�� ���޻(f��2�r�n�+�Yy��$T�<9 �?<$i�0+?��R�U�A�68�B��"׵��������䁬-��ݹ PGz8�S������^[�/1�+aÀ� 37�s$,ݲ��]v���b��=s����Ũ6��$_�L�,�5�$��=mW��"�Xj*�j�%�� ;pe���p�(E��d�'�y�L7�"�I P�e[mu��9r��C"g�徰�X쮻"8���q��#���������#/ޤNR�j"ʪ��4���5�4[�˔��]�N�����
ysv|(BMUԛ%3�U��e�)��P�/��*{�L�Fdz�5�ak�u��NH����M��g��{��Ӆ����K��%�yc�'�_��������g�bHv�GF%�c��6ڇ�׮ �,��*�δ�ɳJYv�s�H����
�VB4�c���_�3��z86���I�{����Qx��m����'���s�n �Q��DW�՞
~���}�Χ�-�����x�↕�M��<�a��Ҭ��.���D�E����`R�X	ՙz�d�F�~c��|{�?o(�&�p�Lx1��[��R�Ay?A�9�@���f��N��{t{��gީ�)�r�0XVv�����P�%%��I*ߑ��l��R��b�@�ir9�iF��.�J�\�/�)�(�H�R끲T�ϟ��G��o�,�YL!��P��ںZs�i���	1�J��s��^@��W�CXS�.ز�X
Vf�x�3Z�����P��T($<h䐪�e�h� / "R]��l����Aajs�w�%�O�Ph豸5��7F�9N+�v#��;{�nU�7�����yF9��҇uUĘ�&�O�4�OD�Ƥ�����׫�>lP�Ȕ���l�E*��b�]��;fXh��k�yA޵LH}��(Ic��D�X+X-��!��G������T��dn]�%)���-��D����P����/N>��f���t9s��e��"�*Gt�?�?<B�V/B���I�+j�yIr�Nu��[Hف���ߘ�:4Cz������!�/.N�:f� ��'��mܨ65P��Uwkrj^Ճ�O�ar����ȋS��v�[�Zj�#q�[�����!��{� z��Y�lo�ے��+�q�VZ$�S�3Ӛ=խ��N���R�"y�^�
�y���{�{BJ�z�Ū@�7�KpU��p��"�?����S4{��C�9wm�~��"è���N���P��%㜰?���B�D������P �粖֜��nhr�q�y�/��0�}܌\h�~�*-uR��3��U�Ӏ�O�R�o���'P��� ��%�S�����^��W�I��TM8��7)삲}$�b�|,nݔ�0'���H��0���Ɠ�8=�0�,8�R�&Z�dN�9_���9G��-���EZ���]5�����=�ُ���kQح�zZ�e�#V4�����'��$��m�ǧ������ B���J\���{��,�+wk �r�ե���T�[t�&k�D�Qy�{t�R����=��7��ӫO�����G��ϪEpć.{wu#~�O9|�e��EvS�����F'�|vI4n��������V]/����&e����ˮ������_#�yON�:��m'.���j�cB�D�����W$G*�^І�Ŷ�-q~l�$�m�2��'d;��\��bΡ�����I��q��(�DΈ<;�ɋ�i�������j��3�l��n �� �C�dr8��Ʋ�x���B����8u�u/��L����y���4�.K�V�~[���c�)Q�����s���V�
�)6a��S���N`8w%��/���a��Kg�y߭HX�XP�@�,�Z����$��ǩ
H$�	YY?�A���&�m�Nx�]1K���E~eq��l����v>�Ĳ2�h��.��t��Z��װY%s�۰"�jQ<��qs���#��+6o��I��]�����H����iI݇`�aҕ��"�\��#Y5��W$��J H��C�nR{�A��vW��R���K}���2���,�f��&B��6�FN9���^��� ��9�$a�2$���A���ɑ�	;wG�B/w��(�
(&l�n@��L}K� �K�%/MC ���{�")�gd2�����7�Cp�W���:jO�t3"�:��8��<c"����� M�����{B86�q�Q��&�"�^�4���d���K7��,0�G)b����g>��\_�];:^SMR�ߍ7z��M9��>{%ꋑY�I泚����6Ǘߠ}u����s�9`~�jR�Hv�-��+���R+���5)���A����d:���:Z,#D��=营��#!�b"*�ɕ�}�K5��q��,Mʈo|J�gnp����ݗc����^xUKyl�%G,?�j�F��S��І���'ֈ���6�Xb&���ԌO�=�(�{&v����[m�9�ZT�#Hq�?@^�U�fG|>�)�$��w���:�=��q�H�/D
��j�UHKd:�nq~��i�?yQ\������(F�;��H��%"H�8fP�%'5�s�����,�\� �]�w|��L�V;��X�Lxz�$X<��!?6w�:�X�l����=-c�S.��ł,F�a{`9�����>�o�Z1y�?vB�^%�W�H�2y���*$�^.x�$�&�S��E��p�b��C���]�����,�oH�%t��2w��T����D�d9~�<g<@R`�S��h�D���]�D����v���H:Č��� W|�d�uC'���/� ��Pe�ܜ�����&K���v[��2�@��4,	���X�?l�We��w��7�1�7�a��ʺdl�9	���Ri$K�:Cb?�*��D\��\1/a@f�S1��Q�E��m�C��W��乧U��0i�㤆B��S�P�pF�3=C.)uei'�V�J���T���� �V���Y s6$���ʶ�2	e�;C߂�qk�ꢚ�X)�g�'�f\XLvnsv��<�A�UuY���i�)��}�0(3�?�G݈��=�� 7�L��g�@��h]����[ Y]Ǐ�SA���I+���=v��y4@�m�����ǥ����y�R�[;��q[7����'��e�tO}c�=�EX����>�,!o���b�I���U����$3p�ۻ
`�v$�S�m��Z�1��1:S�#c,��w ��k�����j��]e�
;q#k�`��ȧV�L['�e��l���T�	VZ�ep3�1s~�w1���� D�c*ٻg|��iG7+�[3,��-*�e���8�J�qvSzǶu1�	K�f��P��-+�Cvf�˛�Un.ze�|�X����7G]�� �|�\�7�a�7���#Dc:��[�q��8��I�O$;$ax�]p�'��qt�d��å����%D� ���:|)T���W�S�r3����R�8��ծ�칸�~�(V�̩p��s}�5<�D��#�
/�03YO��`������Z�"N氧	��BW�^�(5+SJ��cW��4Y�T1"b�;I0c�·K��$�-0�X8�ӈo�S���c(x�!~��v]q����	��d�#��\,�V�����z:�Q��0Ռ��JOĵ%�\�s�;eaT-x�Չ��^����J���_��.���eR��;����%��/�j���JI���L����}IJ����j�N����ʘ�k��I�]�43oImyW|��ё(w�X3��OQoM��V>$��T궳�fЄO�vc��*���l�>����� �IN��3&�V!�ǒ�9N�7�>��f\��]�)
;G`,�)F�Z��^N퍲b����8���@����홦\z@3�X0�P��Z�݇2�[��~Q(B1��0g�����eشk�$����������pm��V�N��N`:��}��S��2Ǝ`�o^riJ\��:�:�K�E��ˋ}i�$=�`�n�7C�ںB��X�Lm<DY׻�Ϡts���z	�3��i%
��K�ڭ��:����w��Z�N}�
�V�6K���Yx��3����wu����y�1�`�z�4E�Bs������D��0iZ'�<���xy̱�TȻ��/�3�*���*����m������r)�i�j�����u�_B<�ݐc����_�y�.��W/.�RI�:q�������`����-�/�V/����|��������_��B��Z;�Pl�Qd�PA�m'�S�R�-0�����{*���Ǻ�L3_��z�����
�gY���Jf�;,��6� ��A��}Ǘ?*�G�'�W�¡^r���� 
�j����9zc����VN_�9f���W	v���B-�����/��[H}"R@����3RÁ���z�W4]�x�&};��nG���P��?y2���R{[ ���Q�|����=ˀ�(b�U�!��� ��Z<]�A�� b��6C�5u��v�R6B̐Y�c�"���U'�rd������%�˦ 8GaHr�1[d�������C���S�$%�eäxY?Ө�1a��?s��S��*"C�#�����p��4��'��Rj����t[)���-B�׽o)k�$�w�Meԙ��s�����TÛ��0lrM��(��y����FG�:���p����I`��r�)z��p�;�x���1}�eջ��b���2~�#@�Uc�_�'Ϯ���w:�/o��`xJ)|�i��^��~�9�)Z�k1ʊ���G����hp�����@����a���� t����b������ݰk�kX�ER���� �d��{����Ҹ��X�;��6�b�ןS%����ԑ�#B2Hm":j@5��y<U^{����� ��gu$G�5����P�E�������+�7�RP�#~Q�p+��Œ&y2��@����d�H��X�N�Yh�ܦZL^�i��@���2�E$�t{��X8Nr�~݀G�I.���g�oH	s��8��BDaA-��/��u��g��J�t��KS�_����9AA����C���Qq;���Ȯc���U��F��qci$;��`�#�()T�Q�fQf1E��ь���K ���\8�o�:@7�Ufh����0S{�W���8��.F!%ՔY�g�VMa��^ǝh�L��OJ�3�b�B*Ӊ��;��r���P�h����bU2����10ےͰ|y��Y@�J~�3�S+���%�0P���]�|�=��r7�lUE���DO�y4Z��?ؒ��z���ڙ��@361KCD�r���J�"||�R�r��Q�|����Ӗ�ݲ���l��S4����׮@��CǶH�����z�	^���HϘ��~~w春q��I�<'��kX놲;���s)՝������������
Rʈ.S4|=b�|>_^��w���Z�v�.}�11P~���o�_�`��?��#G!Cn��U�8�������02rO��$}jj��D�#�h�����L$�I����(�t8������ �%��x���L{�#OOS�'�8M�
|��ɟz� eh-l$bW&�;���rn��{8Lɱ)n"x�툺1�7���㬫�D�I��[P��o*�	�c�d�l�62#S�T`(��iO��#y�5�П��'޿ ��d|x]������,��3c�����j�AKfy��N�s'�NУ5Gu���b���\�D���5�9�Le���6�;`���X��M��x������P'0T�d���yo�;'�`=����sI��r����i�c�LI��K����̋���e�N�h}��}z��,��RJ��޹WON�A�e�9P5P������������ۘ�TՃ��'�ԭH�^���[M�=�lx�7o~����$&�5'�	�`X����m*R�L�	�c��d��D29D����P�F"��{�����de�:F�!�/㰬���$�v��U;�3h��\WN�.(9~
@�y�h)� �ϩ"tE�3�cƥ�6[d.E.4�ClL�.�H�	����l(�wE��12x5����2F�����-Ϫ`���ea�g��&/�=9�j��;E%�T���UU��������`�P�~�ݹr�<��~�k�Kr?m�6h�������z�'��J����t�Y��%{�E�*�네f�#��CYÊ�4�f�W��/X��j�٪�&md�����}�O��HS�Rc�{�@��$���z�V�$��v�B#P�ko��5O� vd�w�~ֿ ��a���,���������B�*zΔՖ��IKO�{��2���|=�e�M}�>�K>� ��z��~7^`#�:�����c$�
��~HT�M���hx\��M_��j>�NRy���c)%�7��D�Ȓb�}�D�W,$ۊ�5˘5KigY�+t�O!�Z3JH<�B(��Ç�?�9dtٍP�ֻ��}I�[\��ڑ`�f.�{`"����fbWz�),_:�uj?M]wz�@��6�ϱ��������$����#� 
Bf[��x��{1��-{��;�{f��jVx�p?��3��w~r��S0�3�r�<��ՙ8�%��y�nYЀ4�!���5�3r�zN�����z��~�G���	0�i�]���Oye���l��И��7��NB1;�FS1��,�C7z��SXa�ǽ��t�K���-��0!�J���~X�A(�$@w5d�2K�e�h6��c!��F��E�v>����_߬��:=C��S��7l��|o���\��X)0���8�Q1c ���ѷ���pܷ���s;Z��<�"��Fg!���1*�'��(?�a�ſzW�xvE��i*<wt���P�w�zԃJ�LH3����-�QC^��T{���k��L�h��ǚ�Y��R@�oD�6!�O��WZ>�I�嬃]h��^��Ǻ~�I�=�5�@���:$��Z� L�B��$|��%+rDŻ��n3��2.��4���x��c��"��N��͢��.��ӟ� ��
H�;J��yc���]:X;;���D]5��P���+m�fUl[���&PI�u$�^��K��+���]h|�Ji)���Ζ�cڿ/E�/������B�V�<���9k�w��o���93p��y�U���x��tn��$!�:Nn�ޡ�.�W5_.Uw̙+���q�P��'<ye��6�Ur��+{��w8*DɽZl1��B�'�ϴ�s�m�y��۠2A�Q�pD2gU�='`�J.Nb�t��-uk�9���{๙��	UE�:���{1<�ňܺ1�_'ǟ/E&�h���X.|�9�W�ʓ�W���x�UZF��l��jy7���~��S�j���T�JpE�<�n�??���o��耵0��������W%B�t}���豦9����"��MW���zjP��`��㤈4 u���M,��w +vM����y�*��I���K�g���MK�������ü�����ҫ_�W�ڂ�u����%@�+�ʞ�_h������d{�A����~��Hz�!\o�E����&7Ff|�u�����Ϲh��5S��Ά��f<�!t��Z���<y����Dz������<� ���,=u=���)2M��X>A�/��F	���e�Ot��{�ub7�/`-�Os�#	Ҁ>�y�n��zV`�tz��ؕ��~qU�ϔPD�zy�3�U��j��fAx��Jbۜ�'�2s���z� �I��!w�3'&��9d�e.np��3r�`_[X׭1p}׸���[+�T�\3�Ց@qxc��ߙu���R����^�@^=S#�N��O����#9�W�J&�i�8���` Ѱ;���y^�aL���C`������቙��.��<P�>�\p+8N��z!_���彜V�4�.�O�zV���a��c�#�㊀�- �4&y�����Ԓ5t|ծ7�aBA�tg�dO����XDU����Oy�w
��	)�8>Lx�Z���3@07���zХ6Ez�[*�u�H�2y�߯;izG�2L�'�W�<�n�hP-M���K[D2�K��Ì�5&�#&0& sP�"ʯ�O���Ɗ`����Z�]v�Ö�p*�+�h�5��6�2�s����p���q2ǁ!������G%�9�������I2���Y����<E�=�m�,�3�a����I��ع�͢X8����ɐ8,�	���3eL�gd���>��~��M�T����Gt{.�Nci���@�mcg�Ð9hYO6+.c�T��X�q���g쏥��-��������c��� ��L���;�u��b�QV��P:���_��i0	M�����}8j2w:�s78�&T�:��)k)�v�"����8 ���:؉Mҙ���/%�!p���V���!!�&bt{h�ŃB�}��&^6f7�ӳ� �X~��c���'L15�35ʈ�gjVW�k����͸Drx�g�D���.Kd��A�d�
,�/P���U���S�6� iNAPæj袼2��z=��^H�t	Qzq~k"%�b��jZ�X��,�h'��i�H1�e�t.��N�#�c!_�|f��ϻS�}�nh�x�R�� ��'��;��#4��ܺ饸�/�Ac-�����	uy��i����!�괱�/ջ=�NcIݯ����=0�Jz�&hq;\���w����U8�W��\@��Ch�ŚDd ���@��W��0x���#��M�o��ݳ���y�!��a�4���@a�a����3�����:���k%��sb3��9ي��>��f��?*��j�6�?6$��v��q�����CW�J�J�Ӊ��>�p	���ڰ�ɟ���K=E�?�h&�F/��=��A�S�ڬ%��Q�ҁ�P%���>�Du�1@i��'�V��'Ѯ��]���I�O�˅��y�[��X�����a�`�,x�����[])�C'*���vR9;����Ғ��O5��g 0:&9!KW1_�HH��b�R��[�
���_����v�k �ڡb��Y�0mѾ"�Z�e�ű� �,:�o}��]k�'l�S��� �ɺ�6�#]l[�}��ȎنQw��V��q��.P��� ��{�MRݽ�R���7\��!GW/b��t����͏h�5��W�?|��A�1��B�B��"���ϑ���`^d E�4,{�*1��_r�!EE�Sk!D ޤB����ӊEu�x��^y�ڍ�*b�w*�H�q�	�џ�>u�i��f �1�%��u���e�"���:��g�Ԅ�e�!(��X|d�����V����=Ƞ�"!5���-)-ކ^�8�3�:�,��`� �A�"qΡ��/o@##�;FCc�s1s(�TZʓ�v)�&XZ��>E|B�f������lF6�������O���լχ�D>�f%(^��t #P�Aʰ �6����Z�w x.I�%���6�Y\�;y���@��$WtRW�b� ����N
��z#�V��sQ��妛<��%�حQ�X)݋���B.�$5�]�{np�����Re�9s�nf#��.�C�א��6��������l�qB�"ʨ���C"!��}��s�
���h�������0�q'5|�`��;,:��zݛ�/ԵS����J��%�$a0X�~�m&W��*y�����T����ߙg�/�$���bB��wr�`���P�>_�:aL���6�}L*�@��0��Q Gz{*]h�~ť�t��{O��T�q�s6�!^��yBGL�"���8�>��<��6�ͮ�w���_��GkeL㢡�m�Ͻ��u�=o1�Z�^��';'}��&i���CT%���� ׮Bq<����y|�xop��z��u2�Ojr;#����� ��^҄��57y�"��l�����}`�v�Ǚ�Tw��������"�&��M�;@l��uf��Z6���|�8v�(��mZw��Q��Φ������z���"������� WK�S&2�>�E]q�Do�L%5ʅ�67�j������i�SQ����*F��p�{(�qSS<?����_,��:lj�U*m�4Y3����:X�6���t��m�-5f�\a�-��8��w�(��zH%�����قk���#�R��,�ldq���
ǣ�|�ق1���&q�/Q�B}Ňb����j��P���z��͹(uu�1��Є_)8��g�S��/5l����)����e�|%�i�����تY���<�Ho��T�1x��W4g%�`y�!cg'b�)xR�:�Ov�FEw���{��{�@m��ϝ��ʤ�x2:�tp�^��_l��� �����d�a����u���6
�H�w�7ؘ�r1��:)�y�
P%�Gq�(!�����*��Y�6Io�E]����
,�~�K�e��&�>�X�ĊmaZ�$��|�0,*$R�$�� ������'��F���v�~m�oo2���/19!mQ���灴�"V(b���iMwg��k 	8�(�ʗ�yg�V�f��nF�Wb����EM����W?p�*�S<��ޟ�o���3$�u����/%�7��
	��}F���߸�q�.����4?U���#X�i�8ժ�}����x)˿\��^��Ɠ���.sܡ��
Gk&�"���o�ָ�H~���P��?նE>Y<���r�S+7`q�6X*mE�{�V��⏛wL�:ֆK|�eD96G�V1"|�]�ͩ��%�ڣ;��#3�������$�r�C�j��
��d�0��<=�C�uz��~=T��zu�h����/rn�6؎�X�܌��z�M5�3`����Ss�>M;{�q�۶���<����L��Ά��իQ4��8�	���fc[�N�|_¯�E�ӛ�G^UP�Z�8�V�O<�OIN�e�I��>�P��.R%�E2L��^��c�l�Fj3����$�~ ��i����})=j��č�Κ��EK�s�ݲ�ѧV �� ����e�tۿ4����-��hW?749 `�O�p:� 7�\W��M$�A|F!�"�o�X��a���W�F6�;E]�+פwъ�k�n��:4�>��f�YM)S䣅W4��.,A��\��G��1�m]A��o�Zu�3~J��ՠp�]}*��Z�������Fr��|�Ӏ4�F���K���o��Z��ۃ�b��  =7q���z�N�,q����]T�N�][�S�����>:,C�q9�6ʒt}�A��1������a����} ��}�ۋ��('�F �)���`�-��$�B�}>�M ����]Y2��K�m��W�.rt�f��:�Pd��6���:r���kgA=���༔�: ����v؇���8��8-�'�|9F�P/��8{�kB:j���A����QJ��E�O�F�x��d|	���?��1W�i,�J��a���B���?��ܷć`ӥXJ�b.��U4�Zjw�-�kZ�e:�HЬ{.y8p�X���!.__�9[����yļ=�����r��]���E2��2`�H��p�/vVcde`F<6 �2�3�K�lk�1��:��h��g.u��tO���D������
A2�D:�Zo�T�w�H�e�0�5r����Sb�k;Hz��f��D���QA�6�\p�C��(�2z3��5��;��Ә�	���ПǮ�� �����Ge�Q!77�*)p�Lܪ�&��d�����I��D�1�� =���Ŭ���m�y��R��I��\�Eb7�8>��>��ޯY��r�q��i}1�^�N�ˍ�0�#�(z��8?���Z8�x�wS(N��oY\A���d^�h� �ҁ�6#��Yd*��d	�S �sa��wF����6ق9 �P.8��w�g	�PȦ�$��{s��u27M@�;��2q�������6�9�[P�]F����Le86:�Ms ]��/���/&YY�?^��4�"(N`��QhCV�(ރgN"��w�o�(��c��5ҋ�;R&���c��Y��i}X�,�����-5=�ĝ:��JDxHj��a���~�}�h~=�:�8�0`�*�x���k{n��k���:7������)}��[���Z����`��*C��z���q��:f����Ղ�#i�Tݯ�����"��=���4N����Β�x�l΋��r@��]��(���l�����Ud5�~���.p�>)	KTt��,��b��}�N��=�:4�������<dU���A��P{?������]D��0Xm�b�5�ĖnQ5�G���>/�*��=Xs��/ H��~�^-F3�L����MO�� �js-LN2��8><�9X����WzCJ���%����ˬH��G�f��f�\B��R�!]�P�x�}�:�LĆ�pB����$����H���ed׃�=
"  u@����ʳ����K�P$:�����#�D�k�e�������[�H�JC? ���9a�����m���a���<�^p~�>7��ѧYJ3����g83�*=�U��MI�S6���c�j�p?�:A��h#P:3.{�<�N�=>]^�+�[eG}�O�PI�%��y��(F�UX��B�MȒE0&O�dS�@�P�h�Xa�rV�щ�AVf��;�[���U�Y���f3�G�n Z��71�����c��Q��h-�E� K0a�ҕ�xn�qr�Ј���m���7V�[`�l2�_eH3�0g�Tw��/�K��I��|����+D L������;Ѹѿ
�����"��x�_N�[l0{���{��K�\t��j@�?�E�uK@�q�Ag6~
̧��i`SO.J2�P0��� Cv5�bKA��*���5g}e�^��1]�nƧ�R[4h��8�p2����L�RJهwl������&>���үk�nYrD��O�9����P��-#�:^'�o�$q%J��w�Jj� k��&�,���<���Ԡ}l�G|P�� �Ԥf��̀�?��zÞA]>��%�ګ�	�B��b�4���#ݝO���ӧAJ�G����;��Ԛ���3�f��} .�۸�[?�J�Ñjfi�������4Ċڬ}��
1Jdg��5}��n!5��'�Sb�*�d�������m%�.�IG�[5��6�� �[�C`3���yΑ�d*�rbWCycur���0g����RFGb�Us ���[�5*WZ>� �f}P��.C�>���#�Y�^�yܦ���!�ɉKt�F��t�����C���-	�
5��_�l�6rຎ�ͷb(���͟��d�ڱ`�rgY!&6�d���^��O?���@Pk3���`#aH��`���)�Aƽ�+U��,K�J=S�Lt���t~�2�E��h&��K���%fR���ܻ�>!9� ��%5$@����v��<vM����6�{���g�A�U��k�I	=�䦯�jt�B�sa3�	|/ď��Qq���2�c��D�dQ���l.ND
?�$P��M��U%\�[(�AW�.3OUhT����B��/<~����
����7��f��H�STi�!&�*l�MC�>_�x��OY�^�Ay Y�g�bb�F�=6�f�l:�Y	f�!4���&�u{ņ�� <��c�b�*���(n�+}�����
����?L>�PuF`ȇ��p� �G���1v0k)1�bZ�T�aӡ´��kX�a�����>�f����ԯf�V�F}��~���C�7�L̈́7%䥒���j�qն%]�X���$����[�؈���	!Jc�����n�W�}���d�~�KM�Z���z9�d�l���+(��t}�1+�M�J'ELM����ӊA_��H_:Ϲ��j.����Ӈ��=d�
dq�,ʙ�2�U(g] ��I�d_[y>�.�97�֍��/U�c�DLwơ�ˡ/!A)߫�#4�i����7�l���&/�E^EAT7s^5TaJ�4�V�P�bb��~ƾ�x��*���S�g_���R#�Uƍ�+�"�1���NL�A���_�Jy�`��#?���4	e��Ėm5������DX}<�R\��!�����tD���/b0����q��ո�/�S,f���z�������\�0�7�@���Ӭ��}�lW��d����໚���p��X�5��mxC�|�`�u�3S�_�͕�L	�e���AT�������UĒ��W��
���U�C8g�Nq�+mµT��X-��=P,E�HJ����iQ41��>a��5�r�ŀ�t	�~�7�,-�W�yC�L���Zbۑ_~��c�
Ml��@��7!�i˴��)K_��(��6kK|�ka!�eLC�z6����.z-H�+�IW�ܰr�3���En��>v���8��6X�sE�Oh��}�C�{�]1�<�M��ѽ�皫����E$�=B�N���������q��Re$,Qk	��*��zƸ�u#TW$��Pz:E�y�<:S�YB�3��F:J�i�^��Y�D|�%���5G�o$��N�_��V�E�T|I����e) X��Wp><�O^�K�+e5&_s�}��'$2�%a�/�Ld�PU���Q�/�Ց���:G�z;s���	ze8�����M���a���XKJ�>��.홟�N���i!�ń�iQD���Sd�t���n���U4:����W��m�q����/�]ٳ��~�ǡ#��pt�}!�i�-6���
�S��?���o|��5*iDc	���n��������9�H�Lo$+�����&^M,�!W��6���������扑0�Q��EF�C+�'�����կ|L�ɧH�]v��(g����hT1?�g�𺸺�ۧVqx"����f:�?�������'���im-t�`�p4��-�P5?�D�e?�y O(?�-�?z�E{x�w���m�U0y�>��9]�dCub�%��Y���pMGֵߵ1�pqsB-=��}��ASi1�ti���a^���P���}9N~���fTov�3�E~�*E�a���hE��I�?���'S�""M=ۯ�0=� C=�슥�� ��4eN�H�Tz񿪉�����+���_�g��4h8�m��00�L^�Lz����	����g���a&0��E�ө	�$�C�����<wS؝�0�\'2�8+�I�0 �ע|/�O6;��DU�����3�2dl����Ri��J�;f��/��1��t%�>B�SP(?��Dc���OiXDMO'JvB]W7-Mq�Z��OD2�l�ڹ�$hT�d=nG'�Xy��ǳ����+�^�uca�i���0����L�_b��/В��v~�P1K���J'���G/�,tuT� ��/���Pxf��4���'���K�����f��������ǵЇ��r�3���l����6�� ^����ˋ~�W�ت���[��ʥ��P���ՍLO���^�TLL�Nw�~T�߽z�R����x{զg�3��{`�;^!x�p%(�	F����� ԋ�<i)�ۻ�uϒܨ�)5��/4�V��/� q���}v�~��5����0�NN���J!=����Td�Mt�i���Ǒ=f��U]���9��ӅWE��1hM#�y4�V�0G�5)����W�/���B�4��-"���S��1Γ��Z��_�]���]ek[:��	��0ԂV؎�4VSk{ҹ[g{d���1� ���/,���i���G��
��|k�&��y�+8��]�����̹��X�9Y�0T�@l�µ�b���2����<�T�!���@��9�Hȁ Gs�$a�o�4Q�"�J��Ny9NQ���xA��$��Ι��4\f�m�c���G��U^��&��p�)�� ��ѧ���HK�p0%���2mwS��K=�*ߏ�*<�k8�&B�!se�t�}�X�&f��nk�`/��׺w��o�C��u%�<�O����P�zc�E��;�|��&;h�Q^a�w,�YE-�hK��`�Y,��B�=\�Bm7y�JN���m�m�n�9��W�;Y_]l�}`�ׂ��^���X�C�;�ŷ;�|\����}��f!ika�Aq~>�O8�KNq��9�*ο �\�SG���JbB������o��󚁟�+7d73z}�����s���!<�֥��&�k	���R��UT�	%X������k������𢫀М �ٵ��ǘ��/�����X�h<�N�ǉ�,��1�z����a�26���ũ�Kcn����v*�yuTO����W��D�i�]Tr�Wo�.~H�YϿ#�HBi����M֐(����J��i%*�Ԩ�S�MV_"?�3es���5f�)����6 �\mL թ;��>\����j�'E�Ҽz�	Hu$��틢�� kp�D	o����k+1X��z��'�>�q]���˭נH�E�$�������I��?8+O���2\�tI�����1������\��9䰨�;�m!O����{�3��D�!�������H����B�� ��B��� �=݉zΫ��A��]c�Iu�o�+P���C������De��A�U�j6HE� 3j�@U91S��%Пj�,��B�]�LZ�/$𨠴��
�U+��$̞���8�P�W$��R �x�[Ͳm����mX1�3/�1 j�<��]��cp0s� ���ױ�;�C��3��j�$?!�p2h�=p�D��|�Bm%�D��u�..0�F�GҮރ@~NXC�� �G~��̱5<���������o�'��`r�x�c\����{(�n�׺��$f3<�p'�Ϙ��g&�_1�Ub�؝E:UR���~	+t.�4�s"���8��\&��J���i�~A�����m�E���;y�ȷ�3�$c�����.I!�������o��;�e.���s���4Ј�z�e�Įa�)Ll�G@����곗/��h�s��Wd�?��z��i���)	�B�LD�G��#+���'��E4��qǍGr:k#�h6����m+�K��1R}�B�MF?iַZ[pA�{���ПDW��0r]TL�wG@�PZv;�O�~RI3;�2㼃�k��R��hiϱZ׶��啑X�\�\d�2�C6�=�P���r����; ��ٿ�8�f<K��C��]E3��]_�;�$u'
{���Q'ԁ�R3�Ȃ�Yg�_3k��h��fs&��֕�η��+�V�y�F��/3��|~�>���=7,&���m��I�b�y�\�@��d�MΨ�Y�R��z��ǚԕĸ��4���j,�.	R�m_�Z)}1��cn}��!/{JQK�>�Q3G9��ilG*;�hD>O����C^_L^��7�|-+����6j���}��+^��HWz**������Ф��nF�J[�V,R1z���f��>j�s�[T�$�h���N��;t_��iJ� �96�I�ڏ�5U�����$�j`}�����P'JǵJL�c��|(" ��х�:���-M�+�>+�ߖ����0<X�� ?�����=��Le�3�z�D�j�4n��g:��8�?Cۥ0��8���>��*�]UV�w(qUű{g�*66�ip��/�:(5��p����!�����u�q�{�&�nNۭЄ�^��k�(`\�*�G�_gr�����f���s2U�����Ƌl��UƳ�
���9��%*�A߮�����u�������E�b�A��8�z���%�`�M�~�WWa'��C)�"#�JJk�O�,�*9U(���	
}�>��]l�ۗ�H��I,A���%�{������>:aq���F'�D��0�BHR.0����N��s��z�$�Ix����>k0ꋹd&��ؙ4���&<w����vm� f�L!q ���w�ȧ�*��|��M	3��݂�DlXTʈ~�������ھ�*.�N��V��M�o��9�:<����� 7�y>��}0@�<)�D��#4_�R�B>4us����\��@��u�N�
w�"�M�8GbA�yV�7�����V���_1���f�Y�y�+Rv�F�A()�g��/�����Cm�i��<�#\밉^�;0������E��[�v�Eg�V=�ƹ*�Q���C��yֿ.<�&0&���ʴزk<U!�1]�Ŧ1O��'�w	��C�e�mg���*G+�2����w�����L�w���Yo�4F��\��g#����(�}7mKK��C�c+~��<_n$�1����w��o����r$���|�k��Om�Iݣ�җ����l�b�&.�%�hJX�F�C"����n�n��x
���k�!��@(����91lz�:\��Ce	���?���]���<��sz��@� ��	�� �Y�ʟ��tM�3-�O}٠��Ӣ�L�f{z֔X=�wr�G�^]���LJ���y(�>9s����њ})0��t[�Xe>k���%�_\�"�X��-ƚFS��{��0��gv�v�t�y�����򆍑�dd�t1iO �l�ܨ��zz���a���ɝ_T̩�|vi���K���8�|��,�f�Y���k��6N��<ND�0�.듟e�T<�3w��Q�|��`?#pX�6�ě�D �R��Sm^*Z�~�kE��$n��� �C���ܠ��Np�k]�u
��2�H�Te���i�ueZ�.��6i�"�hJ�aWo�Cs@�ο��7�A�n����g/��:�/'ٽ��[�"3��A~
_�c^�ܢn0�h�"�ާz ����S�WW��h���Q6~_�)�L��^A�i���Du�p�0a��� ���8�ĻO�ũ�z�L�c~;+�L��ul�=k�ʥ6�,;�2cX/�iC$QY��K��KÆA� ��CQ�����Xq�������_�c��˭g`�:\��v[vh��ǾW����Z\j�0 @� ���Qt��k�������Ua֕[��ط4��?�ń+[B���qsy�ڼ�@�Q�J%��Q��Q)�Z�(�]�,� ��E������¨mߧ�ut�x_$fD��g���(�b�
�]xU�қ�$ TL��C�Ω��|T�}r��Ӳ��֨7���9ᇯ �uA�T�0��-��d�m��a��B�U>)1[9�֕�&v�ZLk1.	Г�?���Ȉ�v�'�8���Т�F��ҟ��dZ�J2d,��y�D�X�Y,^v��s�*���>[g2�{Y��	�c�E$�h�o��y�g�(��H�qߤLQ sw�)O����n$� �-���ø�ҍ�
�\��z���Per�t��v2NJp>�}�T�ϒ�PS�0P�_��Q-D��.`������\W���w����T�}��VTt� /��=
��y2AY��eb��k�so⹃��	�C�{9��"H�F���:��j�]`j�ri=}�B�/���w�Őu�,�l�ؗ�5\�:;\��Zސ��A�Oc�&�c0����gH�I�����sռCv�u�d+Y��~{P��T{A�*E��Ipk	�~=�ޅ��\-Q�2�y>�)�� �z���w�G��ǟl�]��%��������D�M��1`��}՞�X��-�X",�B3Т����)��Ta��=4B��p���'+�*�O��E�����ߥ�.��`��`�RD"~�YPq �"wS��_�$M�~b�צ����Q�$��١)�U䒲��
P1A��,V�W���0��{��f
��~��Yi�;��)�@Xm��튄�(_3ZIo(\�z��Y�Ӥ�RB�&y��dJ�"�,�U�fp<�n�D��L��_#Oi@9$tǛ��ס���s��m�j�S�w����
�H��3��![�f&sA��ݬ+���f'�b1�e��Q�ϚHZ��[�%EZ�a��ӎ��e�K����N�<��J,I��^d�6�nA�T%ER��Ԗ2���r���➝W��y��t̸�Y�#��#/M�_B��)���塈]xL�>Ԉ�3�_z��� �D�3��	�\��*�k8��Ů�������_�&����PAP%�ޜ`~]F���v��Qu#I/bg;�Y�"�kA<�5o�Yo�D�>E( �������[߆����|y���36_�A���0��w�l��[��)4_s�����'(\����_�}G���?#j'�q�m��12?j�k��Q]d�"�'�pI���|��6�1R������>�R��Ӣ(�-PR��E�b�	�~^xu��8�<V�O�l��Et�=�ڟ_U�4��,�Bj�- >p�в���hJ���^������z�Z�L��a�S<2�+{��+=O�P��˹k�=d6��f�e�[��f),� ��j�4���:��I����ѧƠ}�h�]S������$q���1=���1��uE�����ė�8�W�h?��U�#��V�&oT7���j�f0Yë��{غ^v�Q��Z�&"��pG/g+N��PE�[G�<�D�^���@.��$|��$������t+}�QS�T�ب´����u�X�Qz�q���q���7̥�߻��!�ӂ��Ö���H��v��]��ߏ�� Q����ޖ`�y��ih�ǝ��/��x�ՇI�q5�����(2��l�/Mi��1���������$����eޘPv�o�Eg ~�� )n���Z���Г�'�B������>�$�"���ta�SF*ۥZvf��c�[���|�@?zst���=B��
#��>F$\d=\�y���u��f,g�A�K��I_OY��ԩx������
.F�c�Kݡ�NVG�*F_�I�w�0ɻ��2?̝W�Ǵ_�𹻗vW�*�響�R��7�ѻa&j[�Vruu���r!���z�٢��R�@P���i����\��YOo�&:t��E����c��������n�u�xh�wr<C�!��j���Xj���Y��]Ɏ��4f2I��A��m�?�	b������LH����j�	 �zVW�^����\ɧwX����x9����F�m�mz>l�5�>X +B�0w�bI%V\ł�3���}�����T
���2��R�Enw�&)o�Ӽ	K�t�w���%bP
ry���"-�e�A���\�?-_?V�'H���b�����L�גּ!ϲ���de��]�+�"$���>��Z��i[�-w�����]�'-{&n�^�L���<�lk4l�.i�����N�	#b���c0��?�xh��pm�=�4��H*w�9E�T9�L��x4�r_�9���='L�ED�P�:5!��~7^8T�{?�r~�ӄ^`�&�Q&�>C�?ߩU�[�)�G���}~�d�.�0��
`���~D$�w��̘�w�躶&��)���+�����D�]���k�G2���6��d��U̓���E���W���>⢜�;��ڬ�P��=������|���4U� ��q��	�Q6���>1%��)���D/���Rߺ���&)���O��6�og�z�����B��Y������>?7D�
��O�(���s��:�ho=���cJ�2�@�]�Ӕ����D>[��I��xm-:��(�Ba�?b&3���g3�;�b��՞R�kq��_���nN��8�%F���W�[��=D���T3y���_�69������rD���$��JM�%�A�c�4)~��(zcP�WW*��Yl�K�C���4�*��eC͏_�V�*�8�b76�\��r5*T�;�
z+(�8�`K
A�5�Wy��5��^�o�����ns=��8e���7��R�q�8��?+��X���˞���K������|�m������ofZ<Ѻ���8'�dĐ@+.qZ�d~�ٕEE�`a��K���K �͝�q��o��I3�dʉ����%�OM���ʣ`�6�VoG'{�D0#��l�;��������j�^yB6vK
���	f/�M�M�b�5u ��ǈ��}�/	���Wu?ӗ��L'�V���.ů��: _���\t�b�\���&fuᜲ4$�Y��}�~��Xe_�,)�1s5��g�&��#:��k>�^H���9'�p�_�kR'��2��~�7�Ϗ�d�`��
M"��&0w��r>[E��D�Ų��trԡ��`'�u�G��7��]�9�-�9#o����$s)�i �=�	��o>)
��F����^�-E�!��T��Hw�#�N�Fio�y�$�;�r�P7=�ƶT�6��TȭF�$�� �k_�&y!��J���4���I����{<�e��b_C�<ۑ���/�%��S�x'O��y,������b�ޚ��)��ٵ�3�"�HjA�&�I��:{�/�M�/~�K�#Q��V􎍈��1���d����
8P��|$��s4F<,sS�>j
T�A���Oo�0���}<m�pn�	WQ�
�򟔟)��"����+�(������,�@���l46&�um8�L���F[�*K��y ] �(��[BY��vz��h�N�~��srF��?Z(u�p��2�KӍNw^���%�~y���#n`�r)p�6��e��Ų�3���V%�*��(�(���~D2=�=���B�n`v��G���!.�$��|�n����raX4 �|lj�.�V�
@U�Z�n�'c<m����톸��9׀ �~��	�g.##�9�-����������b�},Q�xQϖ#��B/?�~(��S�*�K_�l��yY��0����N,C��/W<�#��D�����wN�iv�?3�DyF����>�;�&��C�SZi9wc�)"��u�4̫�u���J�Y ޛ�%�E���}W�*�o`�Tu^t�_�:ٴ��% g$>.������e8��&�vʷ)יb�4yfI9���g��hUܫ����'8��#��膛w�ۈ�'�v0Z�[U��+���i�������}+Y�boS㕒����ZT��2`v�������!C͝�;������n?�ٶ;"�>u���N���S�Q� ����D���G���č<'���[[3���\�u�ዪ�2!J����<q����������e� X�xe�h�	.c��M��O�
�BT�'vi ���;r�.d�Ƞ�?8���&�Rݍ��2��yUpp�Pq1fo���~�J���ms����}xT�ZH�$�Tl�2�$�wӀ��>�A��$M.I��'sT�y��
6jZ;�=iBe�[���ܸ>���}zG���@��8 Je(�]��-4�ɓ�����h��Đ�͒Y}�{Jd��G�_{?�E�i�C=;��k�^�A��uT���\U�_��6��G�#��k�	4BJBnn�,���zh����}�d���
�8�</�2}�u����8;:�Ta�y]���.J�J���NC��0�rS3��S��R���I���6����&G�an|}<Ŝk�EE[b\������#�x��L�	�(P#��D��ӓ�b�����K�2�j�H>�D��_�h]i���U
-�Q�\o�
8�xX�[���_��!�U�S��`����T�4p�.{��j����?bq��j]�Z��N{���ϲ���>��"��j��H�<M��yy(+�(;�{:���9"I��H��-��&a؉�ӌu@���ѱ_X���Lo����pe�z�T.S0�K��=���yfY��b��;_zC�)}�\~�my>/��Bֻ��ry�>�2_�#ݻv\E�|�y9��F�XM���{�-��xH�#��m���<���d!�Ar����� chJ�/߮%7G�eJ��/L��q�_�8ɼ;��,�v�#D�������.u��:�U�~�kb �e���a����B�_�8�j�"kM����)��h��.�� ��X��6%��z��������VS�`�2)�@@{�g"���J9�Z'����W���E��e:AI۹���Fx�=����Nl��Ԭ���G���#� I��>�j�Ob�MQ����/�F���S��~�i;voy�互lHH�:z��c���o:ңۅ/�+����I�Y���*ھ� ���w�����g�+�d���xB@�B�7�͸�8�<��wFR��;��m�6ȉ�i���wy��Z�o,���Ԕ�Z�!8��/M�M��76_�&�<��+�3;���M͝����#���#��>���w-�k	$�і7$������I���TL���~<�N�f��&�a��C��P�F��K�:#�	��b)?�b71������ �{c7����b������Vu�_�]ڐl5:�	����V�����Hs)n�Rb���F��0/G��Q�q���&뷂�.�D;�r�gqW��:"�|Q��G�@����{A.ьǘ������N?zU������R1o�T[IXu��D�;�'�؋�����)=�s�@�c�"1R�DQn�S5� �y�Z���^PxWS@�O�86}�;�h�@~�T�Z���z����yL"�\�Z�J�2��5�������V$_ˋ��d}í�0�"6V�93�2"n9s~����V�K�(�lx��>b����X@�vvV�#�fN7�K�e�ir-��ªz���o��o���gO���ÚRL�V|��r�-Z���S�ʄ��X�n)�3\{(��P@��Y����G��z�Hu[q-����.�:#`9;��� �ze�jn�R�H��qlx����+t�������l�^�dhr���=K%KA�e�Jё�D����tY��z�c�2mB�5����ֆ-�t<���Şr��ږ�>7��R�@��C�h?00�G�m)�|!��!<Xt��R�.B�&g�k�{WC���c��!D盎��� 1Ӵ��$���Rtd�s8 .^4_R֟�f�����Q�� gs��Ź+ň�==�U��XUP�Y���7y��4Y�o�q�#����]E�C�x�)W�P�ҿ�r=Ga�J���t��m8��9�{���x�����^��夲Ml��JQ|�ի����;��:�2P�z=�)�L&�_�M^�3K1�3���讀tm(�|2= �����I��P4S�6�M ���s�6J�wS<&'�B]@�2�Єug��b���������ༀuJ�T�P��1����*Nj~v�1��C�xP+p-��̐�&�z�dz�e匁��Mxp������8ɢ����-Y��3�-y�gu���9����Ӌ����Ϊs���)�Ecy��lּ�V �j�U�g���&l��X��#v�{��H�/8�b�k�X�63�Km��H7,&��00 ^X�r�˜#i��lm�`��V,w���E�z�0e_N{i�x��,=#��.��z^v��T^.��%�b:���VQ��O1U�b`Xw�<�yI*�+{�fh�;�tn�0Ԝ���9�	���!���knX�C���r5 ���X<X��z�Cx'�� <5���ƶ���Z���a^C�y�^��	W
�|8�~q�#{	g�P�YHS|��O�L�i�X��f�3�xɫf0E�d�a%V�[3Ȯ�d��Q�i/Z9#Gkz���Ww�d�en��B ��������cܡ!-�[���w?������:I�����)+h���cxЏg��C�=2����=	ε�fO�O�6Gt�8JP����_��aU1�0̏���YҺp�7ݔ�sF���/���4a%�|�Z%zg��C�j���n�C��$l�7�)/Y����P��b��`�j� zz�+J�Cu4	|�gF>2�`��\��*��.���Łt��4>�%��/�%��{�-%J�\��!�� ��J�|��g3���)�Uj�-F'v��͵�����u��m���!/t-G����>g��=���6q� ]��C��T���_�p&K�_���a�"���s�O�Mpr.?���u��*����x�P�u�X$$�R+�#��Z���W&���:�1�_'i��h�r�L�|mL[�Iq��G�.�T8t����Q������uV�۔�b(ָ����wM�K,X�-&�K=]��Ʒ,���
���X������6:##� C��%!�w��(��ȸq�6'LTk*�A��c�� �2f�H�g��r�U	�RP��%9�_�Ȭ4��Ͱ�z$�����7~�z����B-B��u�g��=���ËRk�qo*A��l𩧝�aD[�Y�N���Ʀ,q�3����]���"⏖�Uc_}���Bɚ��)�W '9�>��?��Ȥv5W2�w�B�ԃ�!T�qh�׎��=�h+����7����Է�R@Cu���k���%8;E��N�:�)�o+�;�f�(��y�A�m�/]��+� �͞��N�7{xljd�-�+fz� �
���r}���*���V�r��↓������&�����1��s���3��|B���xA��fٍ���*SMA�̡��{1CK�H!���I�ê-�%a��.�
 ����;;2m�=6�G:�����4���i��ۣ��Z�r�3��C�'���dK�N�M���E�NX �]R�p	)�²�?��Ջ/	���0/f�J=��<\)v#�d9)�!{���.�,[�g;a�}�%��Z(�9�bPR��g��5[��n�:�S�*���;�Y���^�����n����P���;}\n�$��ȒxJٵG1�(ԷhCWU��;A��ҞNIDU�:7k��A��6���*�=�e�Hݯs�E�%*0w;�֎��{ӯ�nvuD�����.���"�ZoE�������z(���X�U8[�<,ZS>�Ʊ�=���9s�a���$9���g��kp�v����"$ ١�#�=���#k��'Z�(����U�u�qUY4�{��{�ۏ����T�2����<^��+�%IVm����W�C�@�|AuP���<!I]�*C:E��1'�i�L+��@��,Gȩ�����W؜�0���h<<4�v9�Ei)�g�"@N[���7r��S�v�Q�w�}�ؽ�G�	q`#@���j�Ȱ`��5����#Vhv�paK^bdޏI��Y�?�Q���O���ŹM �����o��J@�5�:�w���St�!�ˌ,=�`���	����*��z�d~6!�,����jm+���(����3zWc	,?ϸ�H@�9�o5���t�o~�Pkv8�Ypӭ���M�̸��_��>G�:L{)Fr?�/b<V�?ש�Hb�*øBm���y7s�1�1��C���6%�(ƺdK��&9�dtr7��]
��@�7EdZW����aM�����ޟ	�7)���H�����J��#]^���K�M�\X�o�5e9
���RD<����nu�܌v�������x~3�F��8�l�Q�{�DT�?�"]=��8
k8Pʀ�z�\�m�����k����a���hn#:u'J�ӻJ��X���J��N��7_���/2�àf��JF :/UZf��H����0�R�_N=̲����m(Mc��{�XKX��i��W�͡9g�p��i��y-o�d9�z�ά�Y;��y1�iLd��ԁ��V�Llq�.���)�-6�-ɜX��0�%1LTm�J�A�2�wB�]�ɧZ���}c�%�9'�r�Ӄ�7^����3[�j��n͛�[�m��q��"�R��x%K�}0l��C���q�Q1<JH���>�iY�~�p���L+n����JXMB�����ʍ�隼���M��S�qH�����Н�ةt����]֤��~y�b��+yȮ��Ȍ%X4�m����N���ju�9q��8'�%?r���K��1�����X�%�HG��=cա���(�\�F��G`�Ա:���[�@��
��6L�!OyS�/<�����z�<W4�|��%��kf�5�(�5��-��}T��	�k5�����;0S�B�pT�&�d$��6p�k���?����c]�i�
ؙ�	<�a�vPn]d�Tc��<L<����'*܌K�(v,o���6����uY�5p}v�!RW	�<������<�j��^is�CS��U�q�#_��7��PX��/_?.����%p�[��+P��nk?ַ�W��y�z��aq����/R���V�{��Ȕ�<��ά�N��L&p�'��Qߑ6�2u'N�\r~Tt�Ĺ��A�>���G9����^Gw�b����u���_�'��z}tY�,�%�����H�Ń���ɶ$��=:$���"i�u:�-zUr 2�D��5���4�I��5�Է��������>��c�?�/�S��I�����/eo�K7�PN������)4Ptu3^���p^�5�Z���eWx���0�1��y�E����
A�����\8���A�`�7Ҿ�-H���4AU��&�v���i6Ӷ&n��.P��'�e�Z,��_��8e1�VI���
� @L���P��]$X�qӔI�Z�#Q,p���J� ��h�+���_�[��&���E-/��3���ZE�D..�E9���8s�vZ�{=o�8�}��1��7Ӭ�� {��t�5��9�Z��@�Rۉ�l�W��j�
.й1gH�Ɂ�k��?�.���h�qrp{�WY�����N7��Ο�[NUQ"`�U<{^0���&\�_�;�<.�QzVOC+&��
..a���
N-�Ŋ�y�k��Ɂ�[�
�	sat�[�҅�< c���a�E�\���<JM>�Y�jl�q 嬦&(�٬�,s�|G�#�.j�R�.�&)�*[�׼`ԯ�>8Ӑ���?�c[@��Hol�|��ycH���C@t���"�6� �)C7�<�l�1�����RYD�����M���p[|u��z��0�O��B���IL'��v=�����*�ߦ�&��[�
L�Ƃ��}
��`�d�zs�p%�2���8�9uS�䥅�.�
>�o�\k�X3^yQ�e}d�G�Ff2�P��fJ���7H�>���K���Ub]ǵل4���������R�Y$K�9vR��D� ��T��ώ����}�	 e��}D@�13Ǻ�r�5mE\塚�w��sN[��˽02B}ސ����g:æP�j#�;A�{���?⠇B�\-��\=%�_���; ��y�.�`��SRr�����.Gֽ�j��ԣ����ɖ�g�5SY43s�΀p88��B��$�����vT���Q���]��Ph�-�SZ��f:�u7��N�\��]�d�� ��f���F�,��s�=WN���@/F���Q���#Y�a�#�ez�-Gw��t�7�u`0X���e�e�n�� d|�7�SS�z�:����f��v��Ο�ɻ�� ��u�'w�X�O^&��(/�R؅���u�k�(C��i߸�X�o4�wJ�79�)��VMm+!׎㆕��� V�2�q�����/�`��2�e!qu���sX��y�H��Zb`���BP.�����������LRq��絛ah:�h�_+�L�u+�:���J�E���5�+M�IߐT�vQ�D���A&6K��R�Q��!���Kt���"j���C��x��YD��6�c*,�Y���{����:�.Ѡ���CG���3j�'au�J�/�Y�_�Ԛ��e�Y�+Z~��lM�%|Ǔ��+��v౿cQ����Y�V��[	�j���������ݬo�!�\�'g�[�I�豘�vPn!���8��'�G����D�wN�C��R�Z ����P�9#����u���96�E_3��H���o݆J��/�`��/�N�S��	�0V
�R���&��k����T(��	T�Qm~��ǉa�2ky��zfBn:�1p~q�&F=�3��^��G�&ZZ>PV�;��ke^��%j%���W���s�V��Kr$�ią9�'2���;{�>��H51���s�E�B�kB�NU�������4��>t��Fr� ���~T�u�`�-��Ձ���E/}w;/�n
��O�*�YE��VU�6�����Ի�<�L������c>�_臀j���ǣ�d�g6�;�Cx7�<=���lۑִ�hTB�{B_�����db?k�Π����F��y	�ORx�@ G�i���'C5�ۨ����?�=�J,3���@HG��>���n��y����Վ���e��Q5:�5a������,�+�Z�t�H�p������Ʈ�(�Dg��Arn���*���\c�w+�/�e���L�#`��c.:s�7��RUhE1�#��������p�����R�i��`�[y�H*5�� â�nG�|w���ѓo����Ew��ٵ�B^�n���@�6����*4_�5�Z�V���b'-������0uV<J�I��M,kO;6��t�5�~���d�L�,"52�M�?v�ㄈו��>N�(O��	��ߧNMY��<��z6���
���oqd!eV��޶#������/�����]����GBn�i��t�ߡ$��q��	8@�|�&E᲻������-u6�V
J����g��XDv����.��Y|�p�o�V#F8z�7T�$��!n�bm%+�&I/p���7ntu�o8���o�V�t�k4��E�u_4��r�G���:���r䭼,#�8�J�w1�pSx��}��>�J�({���Z@w�Yvx� � eD��9�F��S�);�í��d��E^M�2�	��]y=):��P�5OQ�G��Tv?�"�`b�������,���3�	d[(�6�H^y5�\/��e1���*(�����Y`��i�=���(������F]�����?�1�I�� �[���$�Q��<�p��f?��ʡw��Z��TV�0^����{14Y������!	Q�Gʹ���2}O䧖/)=��� Q�-f�d�)��V[��e��X(©U��q���Cy�u���s�>h�%�ػ�s�"��q�;�a�W�;N�����x>K}Sz�1d���<ؠ�'R��D���C�%tp�F�J�޿V,��U�?",PX(�2�� xԜ����Q��1�N�٪�Ƒ��{B�`fw)�v������x��fnǱ�J�]�����FB��n��`8��[���r�qbi�m2�[�*���Q/��s��_*��a�Vj���b���S�M��O���)����{N+r�JDգ:,b|[`䝴�"2�/}XC-F��z��|CJ-t�5��w����J �X�# ,�)�)?i���.5l�\ $�n�E;��Ϣ�U��#������"T���3���k�b��t*@��5�	n�Y<�<�[(����0s���z����S��p-�Y���o���a��0=]x��
���
��6��]L����YI�p�[v�=u��|�D���1��h',�\�ڻ@E69�Ksc�� �Ym���A�cJ/��*@T���1��9�ο�@�>�_��~1���H�?_dj���ѭ���G��28v�P8 +�/=k���\������BA��r:��ɛ�U3��� ��m+ӄX��[��R�b�g�qCi��v�FH������wvځC�S*�&��@G�+�|x}���;ƽ�ߞ�{�T�*nH[a�-Qȍ�jQ��&��$�1�mE��Y���x���@��6���20=��&�>n�f�+��������D�P�����8�#�^a��Ѿ�]�2S­U�4��,p���ƞy�T��4�#�Ǎ��5�#i�~C�4��m4F����7��u8)���I��.�=)=T&(7�o
w2�G�=�O�b��2K�����@���/]O�bB%F>H��Ź)��8�Gb�j����|�h��Ha�mt%�=h�C�4c��oy�S���i�M�5�Њ�_�?����p䃧�[0����e���w����1��/�*�����>�m�'A��O�A������ �$�>�!���k��0�|���l��i�;v�O����:��5;L�ߥv�2msP��+2���5t+��қF��5�h$tI�0Ϋ���Bܷ�.*؀� ���c@k_:�p�V֯�-pM	�i^x wp�4Ԋ4p� qD�uUM��:"��`����
=p������K��C�;6�YC)b5�Ĝ@�7<h%�� ����F"k#�l&�
�R(���=��
��UX.r$�t���؛
�'O��;Bd��Ǎ��Au���!]H�;��JH��@I�ݝf._�0�'<:uT��؋B��%^}��z�^u�.^G}��`�o�>3�34eې�/A06�I����5���3���^7���~���"��:-��I �%�y�b�	�gN��B~^FԖ��;���;aT�/�J�lS7�ʩ�������[�w�"ZjK"}d����N�RfD@�A�?9h��r��&�j�>s�.�4�>!���VA<�gM:����?���>�������&"H��Qig�,i��cmd'S"�ʹ4�<����N����9���k���^���O��ϳ̌���_>8 �G�H��J�����U'#W�E�9	P��H�h�y")�{Xy�i��{�/�*��:�4�"QCUk:Svt����]�<�a�T1 Z'���)��*7�5���� ����;��s�Em��P�����?����/�2�_��R
_�~��)�`� ��	�7N&.�:s�zs	�=�
���Q��Qa���yبi��3 p�+fC�p�"����{��N:�x4����K֑Ԉ�R)bZ�e���H#�0Zכ�c�@�#����{$gi�}��ޭ㰦=��P
mg�է�6\3��@"_��ZW+��e-����z�����dl�oj�w�NS��e�����Y��g-�e@˫�m��":��5�h�m����^���_S��t���g��y��Ng|�~5U��'��a��N���y}Ħ���H"�_#8��A��-�	S\�'WT��K���Y�0��;��h_p��7�Ym�g����Aq�0�۶+�5@�l�a!��t�!=�u�z_�0��I'�l>�L�=�g4�F�@�Q�	��Q��B�	�|�2SI�mk�V��x}2��ȭq���g;���g��'�t6�kL����X�%x�VnT2_������^���C�&�fN٢�q���W�ț���,�#�N!�xf�����W�pXBq�~�f��zU)S�^�}8��yP��V�9�rWWV�=�Ħ�����I(�h" #���d��#T����YK\scH��R�@���J̜8z��>ϕ��:S�D� ��%�t!���Wg�vO�&����I��{�
�I�g,$UݫR�_���5�=J��ܟ���΢ �׮}E���؁�pIo���V(��w����R��^����l�b�T���e�U���NOR��
�e$\풾���4t��Oޱ�H��v�eD�a+��L����om_	��C.A��~�w��V_��YӸ]�6����W��ϧ��lt	\�Y:.=璍	�v%��92��8�)*����7��R=1��T4���5]���=M�B���/l�v�Bw��Ra�/	��i�W�x��â�S��֫��P�j��
cw&C����ٯh���V����Cg�ɆF�y7�߆;��b�X��@��γ",C�\��.�_�qΖv���M����vm��d0�4LWH�ң-=*���zjDG�<^��Rӛ�/!���q�'.���7ш3�&��-��@c��vc��lG͏bQS4�W|�߰���BAHe�knpHNY�[Z`�����3dD(jR
b喬��oɗ���8����Ģ�#
��3ٞG��w�V�Q1���H�M��%���_�Kb����I4��|s7�E�B���j��Avc�᫄��O�6uNx�K�(3t����Y[X�ZW�pm�IUP@�î�?�N�'�g�6�_GC6֍�6\����Xl��ͼR��צ!A^���S���8$�����ӌ�u�ZUu��]a�*e�6,}b-���5M�Gg����f�iR=.�I���H�;s��l�Aĸ�^���Z�����'��\nɳ�Bm�o^6�T[�E&�qu����
�ً#��])���ۗ�M;��u�LH���=�� ���$��#�=�5��^�`	ca�(+pM�L+�.i�.I���Ĩ��?8���G��+;ξG
j���]v����v��.gg�h	I�AY�]S� q*J����r]���M��`��C\SZ@q�|��e��L��e���t�"�#�Dc��Ui�y��$h9���H��,E�>2iŒ.�w�Jޛp��հN��ը-ȍd�T��{��_�8\��n��)��Ο�X��ȵ^�ӌڪK�k�=}O[w�ӕ�G4`��؞O(|~�R4�
c;�<��ȁ���#s0�`�O��`�b)cu�e�'��y��W�*lHe��d�e-�0�+�����F��%_�gQ���#�(�yB���z�G��ְ4,�%��wݱ6�3�����ǈ���Kp7i�	T ��o*�,䮷��� �A���OKܺv֍	����6�2� i�8�ě��6���L)�`�GB�Iq�s�B��ʒ�{mM/�OE��#ԡ�����c���;��mV]�;'�aa�v���:�J�⃆ziY�(�U�ti������ԤX���w67F�i/�ᡗ
�-_Ƹ���1����˺���������Y�Ы��aU��R�ӎa���S���!=+�z���+j�2�I�tN�#�CwP�1E~��"uwaj/h��iG2�3���������amOd�Z��dY�X�o��|�#f�V�����f��u��+%�2�GBg�)��&E�N�iU�U��1���� ȱ�-�|m��QAH��%��M�o�@
�`\�ݞM2k�5����M��G�x�vCK+d+�Z�_���QPZw.-��֑;��?�+�F@��+C���N0���׎^�Y�I�Fn���)w�m%_۾�T`]������짭 ���/������,z��� 1T@����c��b2��x��n�+ٳb�a�����.0gE���g��]��k��؝�u�Zs�8S�82BD���J޼t�>��\�$��ʋc �ci�ÞdArn��	��'w�>���^��o��	_d�)Y��7����pԜ��t׽��Sq8���^��N�4f��C� n��O����!�[5Ӟ�J�����b���͝t���at���ĥ�	�B�h>zf2OR(X����Y�'�r}oYeHɪA��/b���9���5��s?�����g�,K��lL�N��>0F�����3�������؜,p���6������V�Gwpά���L��~bg�B�`�_��	��W6r�����dR�)�%-�@Q�XN�"�9�hm�ߡ�<���Gh|�,�k�|;v�?��.q�鎛|���5�`�6U� �1G���I]A}�h#̈́ZU�д�
����p� ��pY�	V���Hˤ?9���)Q����^u�ɨ�v�gl�P�1|{lP޾�qC�;P�%���Rh���>u��rN���K�$���P�+�*�ʡڝ�C��ҧ	.~,��k���'��<5U9O^�|2_��)3��QO���>��0�V��Q�~5L���E�A8�Pc�v����*���y���@�eucL�av��R�+�pR�,�Md	0 YQ2�>�cL�� #E�m��`��>e���.�=��C�ː~B?�]�����Z�� }1`�q�����I��M��y�|D(Nxz�� ;B�;��� �7Y�.���
���D�=\�x�%v v��Ӎ�9���[����)���x�n��UQ�6p۞��ɠ7�C�~��R6�A���sf�}����6�����#_Oa�O�4�=l"�b��.�
b�ԫ�8�|O�3�����KzQ�PhX�L�����罀����I������f���u�rK�&w"�]@�՘�/\��s'��o�j�M��(�ף)[3?g�e���7�5��T�������4I�����ϵ��
�ϗt��2�ʕ�!Bpe����0�,6��0	k��Y��5�V<��ILF��{��I�EBTO�r
�#�hxS�#i&pѓo\�����9�e<������HOT�d�D��	̺%��\�J��c��}-���8v`L+A��2xk٤�jL�?�n�2v^,���G��8zwB�ă�����?
Yj�	�h5�+=�fz���ĳ�L����w4�'G�4ڵ�*#H�~�(�Igm����\�-G=��`{�O������n�K�{�{�~Q��Ѷ�2�h)HI-��o�§m2c}�s��6���a�t�����6�~Ή�}�v�Q��!���;0	�;����Tg�xV���Q�w�R��1{A���m�7��C�"_x��ۧ_[��0 �r(Dc��ϣ���/]��8:�d��9���a@Ӂ�S1���'�H�Ѕ��O-n\���hR��K���am.ٜ���0�.�y7�&��9���$�%�V|f��	2�\C]9XX��W[�z��r�	����LP"���6n�>��@�M�U;j���mYy�\����ƬJN3	8`Ӂ��-!~l}�j�x��@���K!A�IEL)�Q�)�(iW�g7��aD5��+9�`�K�Kp��6��>�UW
���w����
�M��t����&Ѿ�Cp&��6��`hT0�����_�,nl���mg��phm�S0T�FǟhhɑH��mX�6��{9��z!�����5=ɱ�c֥NAkW�қ�%	A�{����e[dLC�t4hN�i��>\�;ݴ$���		+"Δ����Eo)�
�n�up�c�H3I�p���x�-��a�c�Nr�6�}�S�q�e�x,_��h��B5��I���ؖ!�����S`��ҔS]%��M�hv��K�D�X�E;R���V�*e@�����n��}mU�(P�S���ĭ{m=��1�S'��np��Xy�Yt̲ꢯ�Cܦ�V���YA#n�E����!t�	\#DrK��EA���"�W��u]��<�%���q�O�����=����H� ��]
o�{WZ -�ѿ�.��6��4ԋ9OFE F�ڼ��>�������ʧ� �1:�u�i��	����Fc�.���f6�����c��a���������פ����[t�ti7wxp���J�I�A���\t�8i�"�&FE������8����.e�zEx��c���ڜDbl�ґQ�/`�y��bx�n��q�����Uy�>��5��l�G���xm��Z1-|/������ =����ᡝ37HX%R/U��[�/���y6<%x�\c���I>j�G�}��C���=�Wuu�ǯ����$!��H7�%��mO���;�A��Zk Ӭ� f�#��&�7�* �ڑ�*��͐W��@cVƢp�V����*���=�YNR�H�8ǐ��|� $�0�6�Dǖ��=�aEJ�����T0�ܩ�� �N�v��p�@F��d�B�l\B����9wݱø�KF\�rֲ�6�N�ig0� �c��y��G�!Y��0�;�_�>�y�DEk	�
@K��Gp�Ӳ��(��cZm2N�	��(#Ԭ��&Q�SH��"���묎��9#��`�B��.�h3z<(uq�T_*9/	��X+=������N�DM�jd��cʓ(�Lv���'��>4��ϝC k�ʑ�0I��)�D�H���{`Ci��q%���������{����`��d .Lh�c}gB<����<b�
��'�s;�ON��$��X/��O|t�S�i�"�%�ä��'�������OȼJ�͖���c՚IJ(d��y� �oΜ�C�؀.��fB^:�z����w�wJ�B$�&s]��G�7F�u��Nf1���� ��?)�n/�'V��t�_S�SC���qv�T��1_�+�����?zxc�3_m����!��\Q�:K����	OT��a�g�Ăj�������LXeb	r9���f�3~G�FZ��
��,83�/=���2K~}ω,�Qk^k���-=㬅4���q���Z��6��}9
�Y�u��7�r�*��.DpK��բ�7@=XdB{;X0kژ���)7� ��?:m����/RSR�����q��w�> 5�v\R��gW� �2+^Y��s����ĈC�(�o3��L ب[cXPgQqkg��4�©ߨ��"�z%�ɰ�b&rճ��{��(v3�Q[�>��7l���8��Q���N��T��_����6���]���E˯T"��@W��~{^���������sjQt�p�ۛk�J�M�⮏�򍬒Z���%��U��	�Y�]��5K�33�`�Ժp{�B5#�aJ���e��j�p|\�u����v&0��=Δ���8̮t��]�s�HK��W���O���Y]��Oy'?��	y~�cy)�g�iH-=Ll�tP�@�&�ԕ`�D��z��=�2�9��s�b@�W�G���X蟛���0����CH�;*P@�=����DE+�'�/�p�[LM�hiji%���TJM�q6��n+S-�Pc{�����@��6U+�]��뇥܂�7)3���Uja�-Dn�m�ko���8<Ug��lW�����z�D 4�{���(Nj7_� U�O _�	~��ik�/m�Cb�7`B,�~��M+��v�QO���Ԟڽ��_K�8�F�/��eM�ht	�!g��.�N_�)��IF�Yd�z�al��oe�B�z�K��A~lTL�TN��f[�v!�?�[N<
8T��m5u:eޚJ0E�R�-�똴��F�]!���jC)W��,�/'����_op�����>���i���(H�W��k����b�Y����5�1�l�:-,p:�x�'D��4�����i�o玢=\��;�� .,ۋ{I4 ����8.U�=Uhٻ�B}p9�
���1������s��2ƙ2[����|��uԄ�q��>��3�M�]����0���엟~�7U�M�C5H���iQ�g�,���;�P�2Q�ʭ&~�qR�=��F3�pY���4y\��
,���tkH��c�*��~�3WV[ZN�����iq����7�e�59X� s���u����G,(sp�� ���=�bC�� �H}\D����̼8p�`� �(m�m�|}��BC9uz~�9̗̎��<�@�w&��U��.���:k��ܓ���q3	�\�"�1�r5��r&td~=*�F��B��B�pY����%��`Za��!^TZ����c��S�%#�ͦ�C�0�n�����u��0��u9�A���Ȕ��M)qUf7A��]2{;8�1B�Ga�A�ヤ�룹�by� �(ᄄ5{�/jv��!/����{	�^gC9��iW�$&;[e���n�IJm� �3�j�V8x�F�c.���q5��;ژ�9��wf�2̮�-1�E�/���yj��(�m��|��]��M9�N�ӌ�|�����8�m�������_3﫟i���W���Q�_�����Z6�+���Z~�R�^l�,=�^��*Yc�~�����/yi��d���&#b��l[�o��EG�90?���u�pM��",N��!����jJ���wv���$���B�o\&�L%�ū�����K��#U����� u��:��R�M��?�t�@I��<�Ze]�@t*�T��X
eԷuŽ
#�m�ٴȺ0�Fڛ<xO�u����`��,@���!A��_�ޟ�����3,��>�FPǰ��(���7s��,]9�1Ł75�B���
�Z�ˌ;�H&rE����:ݎj��C����Ԟ&֫�vW-�aNI���.�U�����H��B�}5���W��s{����>|R������;��/�0�i��]���=�{�wC��/?�}(���L�يb�+l�=�7�
i\�E�N��I$,��>��5�R�u�	y�/�����N9==�����-	.H���<���� ��M�#�l�m��| ʝO�+���Z(g��s7�g�]cM��� �政��~b��Q�j�����pF�@ؗ�������Z��\G=���h�I�ܜu�&}P���$��rT1���B���h�z�ޛ$T�� �k�&1�����g�;�Á����i��ٍ������	ϣ5J�k����O��b�����q�(ʚhu�-�
0��U(�����槣�<�r�>��2���U|K��x�"���;�h<d��^dv�´D/�q�g�,]�����v�Q��j�e�������m�}y��BSq��C"�ҹi���4�	��o�"h��7���ÑjN�$���0��d�@�s	���AD}�T:���U#�����u[�f��	��ZƉ�H��e&��<�Ar�g��g[�V�����Z��P��7uu�*(��#� �?Pj�~��{��("�}S���醴ǆ%ii���{�Zn�#��_H�N�ƽH�K����뺱���ApD���T
�W�zcVUg�����(�>�����ɏp$�ire�oz����S�{��	!4x�+xZ���2I�y�8�O��*ܗ��%d��D�B!����Ж��
^���ҧ����l�2V��喡��	G�g~Ļ.3lD,�F�~L�V��F";���O���_:`�P��4���2����DM:鴺�Z���Z��c<(/q_N�@�% �2
�!"��bg:c2�M ��N|���0ϾĬyf9�qfs���*~���wq����,U�����Ň9�$|*|Y[���f����ksrz���0�����an��;[�l�&�Yc>��@��<��R� N�E�h��e'��Y+u��
>vU3:�rk��lC_C-�RI�9��?qN�%��9`h�0I�}*j�T�9F��Í��̯&��}��Ej"\�[�_迡}�$<������<}q�^,Y�'I
���J��{_mX��-�A���D���b�����	)���d������kWtȋ�.��u��K��+�*} �������kU{��M^��Ga@;?b�O6�O&#,����w!�^��qV�k�裠�����0s�oM0� �qi��1S��g@�R!U��Ԍ�\�Cl��>�C����~���� 6��� c%[��̉��ni��(V+Y����=�!M?�����f�T�?�3�ѓ$-�%b0���s	��iq���������#a���Һ<7�B5N8� F�v���#'b!ˉ�8��/�y1u˙�Vf��n$�7Bel���/.�yA^����ۘ>.�^���Մ�b:C?%�%w(��ϛ����:�r�h�����o|���"���%U��}��tw�z�>3ճ��.�yA�s��Y@tr!ng�x�XjT����-Fd�s�u�y��i!,ci�7R� ��Ѓ����9O�Y��h� ����O欠����^-KUgx���lA%ߛݿ� f� v�� G��c	�ȁr�sT��0ޟ�ש�����̓Je��\�o�y/��R������Q�,.	�}ߘ����)�tU���}��6A�Sv��k�觡-00
�2)�^'�\ �lV���CCcW)�6X���a���ZC����]�U�Д��� D��y�&���l�Z�S>����w�s�$�H�T�_�Um�e�)�ʛ�M��O�]�� �7(Q�������<��C)Z"rz�e�V}1�Q��(�i�>-̄��4��76��m���w&%|Fx��&��0D�[�Z#��$N�"(,/(�*�*���e&�����,��?�iB��/�\����fo�B��k�NtlDi�opx�? �3���X�IByw�K�~9�����y�C��u�#�NQ��,Y�	f�]��,=O;|�|� ��;b�W��iN/�+.����7�9�% &���H��`K#$Zz��U�b�TF�I�g�Қ����.M`�ʩ�Z(��&��S؍�
p�qf��n�H�K��mw��b�ƚ%�n��l�w�2.rl��6�T7�P>p"�G^!� ����b3M{sx�.uZ�g��cϿ�9��Zt" ����m�d�޵A�,�V���l�R�bUq|0�wFf��)>�$i��L����,�*��b,�6!vSZI��Z�a�����;\�y�'���6�I�JG����6��U�؀ghh�sQH�l`lV��e �z"��XM
��y�ھE�[���$я�K'.��_�E(�V�M�Cz4?�٦���$����יr�������&��n����tJ����Ҷ��js'9�[ZE�U��68���wlJu�|(.nLh�*׌�(�^�ӛD6r�i����Xu�Ő���>u'HK7>�0��M&�e�q'�\���9<��Ƙ>��@%��^����S�m�t��%�Z5N�qF�n+�_d��$UI^a��������Zܻ�f���&]g�0,�C<�C���d��T��`:��"��N�賘�o�w=𷶯��jѸ��3-5-���7���TV=hY�$��l-k�}x*{��?|�$ރ� ��+��S|PA�S1b/>������r�'&c�T�NJ�:�@x(6~iU�6Z��,O���?������M >�0pl|�������D['�R\�Q����Ȯ�j��n�h�3�,4�*~����m�5Q��%L-I^o��˾��$1C�\K����5�:['l�;7`s��b�t�;��U�gh��_����םF���K���s#����#.Dj��G9D֪��_*�L��P^ �o ʛЌ� ����Y��$b��V�	����yett���R�:���Q�h��Ϥ�h����L|)��U!]�a�f��b�Gv_Y`w�t���<��������(#�"��	$+�*ͱ����a����y��$�|���ʛ������P� ������@(�M��&���:���)�j��m(C����K!b�<*L�����m䞋�"�^M*r���}�>�,��?/�]���A�m�٫^�n}���2��<���7����>�`R֖���{�������ࡂi��� �cN��mAP%��_���HE�׉-�m���^(ɣ��d�y巃�LF�[��h��o����j���c�U�I�p��K�;�ǇA��<kD`ٷv{!y�V2�)@�՛�bՌ�X,�� (>�O���l�I"V��G�0{�s�{�H+��z|PK�5`��Mhg!����j�DN bY6���%aآ�v��B��!uч�~s ��l�vp�z?����OK�%&rȲ[�g_���S��&
������x�py��o!������0,�@�7-���'8�iTQ2s��$F2�6`M��Z����\Rl"�E�HH4��0؁?�ϚQ4G� fF<� ��ٺ�D��2f	]����-�Y�j��=��Eu���M�D����s� ���5�zo��#�*;�����D�
(Ҁb��1�����G`�U|���h�$)��>�P���N6��'����r��#Aj� V0#����id�l�l��J���r�,D�.���BĆ�Jh�͚�N����Y"f�J/�I2�	�V��枸%��>�"�w�Е}��Dv�Q�ٯ���@a����JFi��>�be 5�M&'���W�\�H�!�����_@/�&Y��X���p?���'g]���������s	K��iI.']���Rr>8�r�*�������PL'��'�וf[�J��pd�c+0-�Ǣa�}
��-a�{S�(JV�Bg��9r?�=�q��$�QM.2^H8��S�+-���"z�%�����)��m6��P�x�����3���'E{��m6�%��������v�҆�	8$e�{@ɐlg��X��,i���g�#��$��{*%�Է����<0�b2�͔�aiR~��{� (�˫v��I��j$iy��3T�2�Ov{:�Rհ����2D�[�Y*K2ߔA���U�N�tK�L1A��0��f�(� KN5c�_FU�j�=O@��It���3c�I<�2P�LV
m�ǩ)�92�Iʼw�d���#Z*��O�jƏ�8`�uV�g����.1^���J��?q�!�i�d��us�����؆g�D�|$]���K T�
�Y���ݸJ>':"}c3�`�)Ҝ����`EJ��4c$GP�*�T��*E����r.M�+�N���� �j�-ty���.'��@���fsJ��s,��%��ₗ����nJ��~آ7+BM]���X�'}�:O��ƻ�7F�5�`�Ӱ[[<#%�j��e�\X*a����rb���Ah�����M�L�4kϛѸ\����h�#C$X�By��8-��I�v�E��o:�	�-�H��)G]�E
<(�(~�x�?w��29�3czg+OI:=�_����i$�hq�|�D�S7t����QW娩���{��#�j�⌷�� o�?}.�����I@L�9E�����H��"���녏����Dm���b�S�(�C_�W����oZ2��ǐc����v}3wf�T�@�]'�_�����i�#�7�$�>1!���zn��5���A���.�2L�	Ȝ/�x�X�:0�u��<yƕ��ȉ}�N�B��X �&(G4�ur� )������Y�No�{�&��-�
���y�'C�e���i7N���|zpO�l�-S��q��B`b9���ľ�����v"�:��nA|D�J$���	��`�*W���_s�=�6I�1����71�d@��祇uڗ�jɍe�eG��a�
O���2;S��e� +'b��=��R�G?k?�=��%�]�s}�9zm�:�b���c�^���?����RLXe-�CC��*��Db�疟.���+7�>�b�A!��K"	�nk<1ɴmhe���}z^&������d��p'���8Q'ű8)4j��	�y݇�ۧK��oEF������6��l���p���w�󈛀�4�w�B�=�Dc!���[�����92�7����$�W"�C���t�&���*q��G�)$Puӣ�juXϹ2�?�iCV���_�|������F}�7�%�j��k�^�G��.;9�=���e%��e�#g�Q�{Qd(�K1�|5�.[�� 1@���^�J�O��k�ᕅ�����d�* LO�ms��\C�y*_:����u��q%��(��6�dR���c���}e�"�����%cRV�048�o�"������{��cɱ�2��{����"�(�3ߕ�"<�hD�"�b�������Ғ(7�F�ӱ�]}�uVY�`�7���sK�j;>F���s�뤸�P�5h�7����,D�㳸We�}���R������(�s�A��V��d�.kr8��I4���Ɖ��z~A�jH����N���b��J�g!�x�&�er!`ʇ�e�������4�5Sq��5��Fk�������	�N�b��3*�2ZM2r��Lf$������ɹ�,�peW�fx��&�/���h�0����n�M$��E$�1
O@?���-�����g�'My{MVv�Q<���
�� Ω�3��#_ -7����s9N��vK��݈H�z"�Q2����p~4}-N�ΙN������[�S��Ԗ��u���u-�މ�!�N���b2\X��ϼ�dպ�!�K����3?��%]�2�r�}w�Ⱦ/�hs��m2�<F7*Cw�Z�DN�_+gsb
��?Dt��O���z�"��8_'5Ns�[H�#���ٓ8Vi��Ib����4����v$<^�0nC���L�~}����B���-���Цak��_�lK���1�	vz�S���z��K���Q6���1s�Q�b`��gi$�L�^�vs��pNߘsd~ᙷ"��z ��L7}A�"�Y�\c	��[�b���V1ij�8�(L�����oR)I��qK=���q�+��>9��V��|���}&ĕYUe%(�h5����Ka�<K�@�(�nJ]�<��E$\�nW�Q�����đ������*M
?�_��������[�C-)�`��c�qN�d����� V'���g@s�N�B^�!�����g��춂	�/���ҋ���P�^�Y;CB�d>hF��3�ˠ�� 4�����<��,_�?1���f-��7K1����K��h���Z�r�D��q�4�x�CA�e��f#0Y_A�7;R�$�{lE��j���O����K+�M_(nrKyލ㑄�3项��(��4[���֯!u����M��0�� U��>����4�/����u#�+*έ�=�\�[�.�d���7l����t�c��^�F�h�C˶R�<���y�$���</�yc�CN���Жʯ��t��W��Ij#�o��=0ˁ�OGYO�0�涆�t�)��Y�ٚ�)��j���x>���9���QU�5:0���B]��.�X2�~�K�:��UZ;=��w����A�ʒ4�3%�m����,n/���`y�m�_#�B��������'X��>��yغSe'�#��Q���2%uZ���3�I��<n�N����^4&���Qp�	<̎�� 5�T�����H,ͱԗ�q���#v=��N����x�g�J��c]C�.����>��X���tu�>p �cw�rǶr��>�ɅV���T> ���>����N6��t�Н�И���'��Zn�<� ��F^���$���q���u���������t�.TZ�U�fc�dƸ02T�^�' �}���P����z��%��-�WA��8�2Ev�O���mN���i��V��p������%A���k�`��K�}>�/~6�9\��0-=_rי�� G�
�'�w��P�Ix�1E0n��b���XEѕHTRU�En���m`�l�ۘ6��3�
������@�v�3�	g���ܐ���06Mtc0�&S<�vS�~̬q��%Rv��
5>�n���v���G��δ��b�K�����Bۿ�GS.�%�A_X���G�<����16�b��f,d�����<	���\�T��i���N���2w����i�伀�ATO!jC�:�][����B��D|md-�Wo�vꁡ�>Z�m�q@fI^bg�#r��+R��&�:�B��҂�4�{��DO�ܼ��&���Ig�r��q@�U���g�p �b�܆0�h�\ȋE��=�G���X�[SVlc���$�R�lc?�8��ʃۄv
�b��];���|�GPS�jBU��g�6a��!�y���!����JdPmY�[��T,O���Ι�f������g��8!IHP����&t�#��x���kRP��i�� S-^Lc�T���?��x"��lG!a�T��u�E,,2���0��rhͫ�,�7�=5Uf-켻E���#�V00��&��.u���RvA��ug5R�����Pz/X�ЕH�;�����]�5�?��-���Z�6�p٧r�@Dw�[�������@�{�U��,�MT��;P�h���ʹ�#�0k��Ŷ;}�W��W�y��<�"�iH���+��K���]�k���D��+���=�x?�Edqi9y$-�>P�  O��8�v�*?�H�X���=JI`���h�l��2��Z�		��ޤzb=��|w�ɶK^>җ\juka ��������lxz  ��l�C��>v��/���h��lP��^���H3�d:R}�<�OE�|��ZԼ����"�=��h_��'5*��4�<���o����ubI�2��jj^�_ђt��׭�Ё��.GY�.��I��}��)�#è�게sڅ���e���)2s�f���&�S�f�=v> �g�/� Fs�!2O�*�5~�:D����WQ�&5!��Y�l��XN	�a����T�NP�/x�9�洬��	,��t�m�꽪�j��ru�ݐQ^�4��%!���������)e X*�� ^��?Alvn�8V�=�^��8��?�B�zz=쿒GT6�=ZDhc�
�)nZ���}X��%[]O_X^:����g�^Z��.5<6Ќ��9� �z���w�{uf w��A�fiG�"�ݙ�* �}����<4o�6���\��܇�Zkkˠ����9�\�>bD{�����Rs���Us���n����:ν��~w�2E����{`��_�lȃ���>x�&�jd��1� �S@�^v$#o|��1 ~i����A�=������f�NR���eyk�� r�p�T�� 9�y���5Ķs9Q��>ɝ)��FA��2�(��}��g���Į�"�R�5�	���nZ��|� ���A���! �y�@0�T"g��'�	�J�F`q���R,����s�,,k�NG�_tb���h%�����E��֯�#u��"�(y�\��,H9�̌ �;PR �l�	��=�?<�b�l�.�?�t���ջ�J�?,���p@(�brCA��L���BCE��a�Z���p�~א#S9H��6Q=P��D_�аw�����f�{:�*�4p��wID���t?����;�Ӭ��4�Br5�� �tAu�9���!��u�t�=K�ԣ7�|��Z�?�3�4NK8��z��[15ZP��"b�HՑ�Ȁi�f�S�/<x���XXF�E�K�WXa���b!��f~�_
�U����1	��P=dF���9i0<�����0�8D�5��eˈ�af�|�̛��F\�0K��!�ѨH�Y�7Ҙ���$c%0)��G	J<3�j^��wc��u:0�ir�ڦ�/�DΧ��XŞ�x����M{�V�>�q������n�K��7��FD�2c��f�R�RI�oU�=̙c;l��I�^P�Lv�3��[�t���U`�Q��	����Ϯ.��&��\C9B��Hb\����(_�eӛ%��?�R���!+��RC�цA߈��b_.���+	�ܑ�T���ԡG}{n������A�����"�,�W��Z7^3��"������)��n��}�)
D}<��I��3�"�g��M�b<{^�]K����_'����Tb�����xjuV�!��ײ���H#�-�rc�Da{uB�X��q����?B͐C�'c�=�'6z�I��{�P?Jr����
���Olɡ+����3&�5l�<^*�'���ޣQe��w�ױ�
��1�Po<F%���X@Cl���T�vEa�*�ᕾ�?��xFp����5$,�A��L��!8pg/u��ڬَ�%q��k�{4kFY�,�}�f����A����.�p~��[�3.IQW�y`�S�[~]+�H���Ŀhe`���Wel�ʊF�!2�fT�v��U"a~.K��Do`*����G����U�m�X
�A�p.�6�:��CǬ߬��\[����!<e�]���Zm�b��Up70crȶ�h���Rq�@����1��q� @�M����	�[�l�P��Y�F��mb̠(�Å�h;{"Bz
�1��}��YgR�L�a��4@������F�p)����Ϊ�)ܒSr���q�9�m��G�q)e (kv3�5�C$~�:k�,���,tI�;��B��V���K�L���x���bC�A���p�V�aubz��h���5^��bp���9^0�Nۣ�{��Ӊ�4��Ԉ·�P^���ゲQYx�(���%�nr�Q���˵&�޺�V�����9D�Jeyb-��S���o�ep��ǻak�28�|̸z��T4(���t�O��h�
7`�����IPzޡ��x���=a�Qu���Ԑ%v��d� 9�**�od �=��B�1��R |�]&�of'd9��I�/��|�F��v�Çޑ	A~?�h������^Q���Ho�a��wSZ�WH��>�C%�V�,[��T��9-�A�TZK(� ��Ee�W�CZk�݁�����d��X�pq�j��"-qW8^R�)Lr�V?Ё�	�ȃ-����h uϹ�(��	2��"�Hm((y����k��4�����L���b��F4���ZF3�wҩr?R:cc�#5�UdB	5g.�j� �Z�%j���I9w�ݭ��O�Q�o�=7�"�����CŢ���@�����G=N s�D��_&ŃuQ���i��"��=ǿ�(|���"L�=��x}^Q�$��T=� a+K��B�wH|�(��M�����Z&�,)�7]d#�dˇ��Ϙ�$<U�G���}������I��4�h[Z<�8��H�`fCZ��J�h���(���M��(|/��v��Z�,\����r �[Nt���ʹ���9e����ͦ��b����E/�h<�V(!H	�ڪ���85�m� ��}	�R(%$����6������^
�E�8L�[��.rM��`M�\0n�1����'��L� ���H���m�����y�"���=ɜ��9�;E �ek��ޗ���?:���nGy���U�0�*�e%�����\~jhV�.v�i�Q��~�c�m��$\n�,��d�d%���c��#�� 1� ǝ{�����$�aK_�n�_#�|:���W��C���{�*O����8to�����p��_����FP�K�H��솫l[�[1n�\�iF��_�ɇG��%�2��<]�g�J��g�и�6��"�]��U�$�=�?a`yN���.=�d8��K~�3�#�)Q��@����f�!��:��"7�������p ��u]����Q�����[�����x��cd�`�d���o��?��<���U�N@��>^n���飊æ�m�y��/n�Wu橳��=;�F�Aݼ @�����-�ؑ���Ư��P������C/wB���n�lZGdi��B����D:��՟wۤ��Z����)h�<�9���T$��u���9.��z�u;����r�y���XUl:��L�4=9�]����)���qY���S&�Z���������r��!��>AaO�(�P8QL���&c-�s���\d;�ޗB�:S�]s�`�j���~g�x�D�/���5pM�\�&E�r Fs�!��A�TSv�d��9�2(n��� �g�b�n����\��]�+��ۆ����ER�S� ��tc���CN���*���p�OZXFܙ5�hu�uS��捏J��;L-I{��=G�Z2��Cr���6y� ��#U�	��C���?'�S���0�Ե��)���a]��*�]_`��܋C��.���P�A( �(L .T��?�w�C�M3��L(��b/΂r�Vɧ[Ҷv<~B��zR�F��n�$��?WV������]�<������o��<I�V�I+_�$>Q6Dح���e��680������`<	�$ú��)
f^�,�z�H�7btd�f:	d�d��� z����~�%i��?I�9M
%��4n)�&���ԻD��9p/1A�=�k�F����I,���m��\�T6�~ј�H����f�6i�P@������5D�{S��q��+�;g� �p��jL5�Vawjm]���Ea����{&��DL�_̒� ��W��,6���A,�������}!�#�c�:�M�:��'��V� 5�M[����2�������Z��@8C�1.����`�zӓ���a
�Wtf+ЌZ������%u2Ÿ*���U��S�X�o��ڀ��SUh{.�-L�3&R(�چ$�+� 6��CG�^ֿ�v�%21 �Alq��
�4z�	ۤ[�wyp��XF���,W�ew��͠`�X�/��M��'0��0A%b�"p��	 ��lÄc;����6�	oX~)�����J�3Q:H"��*
Ħ�z������A��S+{(��7�ߜ��[���'8HK�;Y�m��gkL	%�x2 ���;��S�R��&��^�F!�x5��P^U��[ԩIHaH�VN�Xh�S����60��	��_�j�N;'��jg�(�P�f��YK��jX��zs�C'��*�w�ۖ�x�����M��w�K�= q싢�75�R��h��%�U���b{˪�^�;����걉�����rV�4}ۜ����d ׄ�.GR�8�}so��WΞёu$bZ=��- ф��\��߇2��]2�G��"{¼�kP~X��f!��~L�О�!Ih%!�Rg7���%&�yG6�:�;<�f?�4�Rp'�x~��b)ճ�9�#+���"g4[��˭y+���6Z�4��g�2HJ82Ǌ"�pq&'��%yRy��wm]%�P�:�
�dV �kZ�t4ט/.����԰Y;�z�c�$<Sն�,^��%��}����֦�栺�0��ԁ���'%mf�cc��3fzc��K4c�7xc��=�Z1��������#���
�����2l��".\����wӥ:L��7�q'ݘm����hP����-!��\����73:^ڙ�F�a� _��aӬ�frD�7zf.�ή��'�1F{-ؒ��2GS֮o�c�����f�XV�}>vD�[�!��B�`H=zy̼�i�5љ�.�����<�zL��v3-�\��d�=ha=i����t�%��6����˼0��ґ�|�"S�[�+I��4��1��m���H%>$?��fg�]/���_�����\��1b�����[X��fn&���Fvp�z^an�����#|��"�R��)�ڟ�.	o����6����|���(�ݫӃ��OJ�Ù�54� W�����i{���i�nǎq�%���^9;T'Ѯ_����S��?MjA"X����+���)��8����ۊ��Jؐ
�׽�$�\��BU���5��	O�/e5H��4�E�V g�/�?�z{����BaUʖ�]�sܫJ;/ �7d�&���p�=ıj�t[}M�'�y�O��R ��Eh(�>���u�G;��z@D�3�)�z��cs$�P^{:���n���ѐ��j��>��{m+�#Uc2f���E��_��n�J10Cw�2���Ǐqq<���3�ڿl~#��� Bo�S�d%�«��:��a|���Rb�,p�R8�v������u+Lh�u�㮠���ql"_0 1����B	D�M��b#O�u��m�����K-tL�ߞ :��M���v_"���S}i�}�S0;}%_Gl�ڽ]������-�c�O��!��M��:%�d�a����0`ң�B�c��aY�x�ڤy����P���%�M2P���c�B��U��/���o�}K�N^�|#����J:k4��vs�kLˢ&Ι�7ݞ~��̀�Ң�aNn�@)9�W�;�������l�`o):�_Ç�a�Iw���,*�,��1;�W\Xp�AX,�H������h��Cv�� ���CK����S�@��ٌ�.m�ǜip���ц%���dɧZ�I��8'��dc_t��F��@��f�Z�ޞ������#ŎoDϪ�*UL��"�I���Ax�DMy;�qq#���75�U���Q�#T�w[̅�fm��1/�U�{��W �Z�v��o����`O�þ�UM.��(�8e;)7nխ��R-1�@3��Z����zO^2���V,�ˍ���6?T���?����Jֽ_�������G�XRoY@���|Ws؄�-��Xڢ�eT8	��Ia�T45��� pS����%�3M�c[��/����G��=�7�v�29A�Ū�Bcd�����0p\^[�U��hg�@K���MG<���f�Ti�kFܑ:�	�GS�+	1���9��-R�n#���,��ε�|Ă���8���8?!��w=�e�n��Fxs���Q2�m�2
jz��z���a�D4�����?��Yi��W��ٞԺ�e�0B�������Z'��u�0Ek�^�<�n�دQ5��Nx2�@�~ⰰ�~�2���VҴ]"5���"{�d���j�y���CSx�>�0�Suw���G܌�Z)����k�Q$P�ߠ�4K��'����D�+*]δ�Q7������iu�,��{����*�5j���Z�]��Г)8�O2�w�-8g�k-�B�U���.�����2����(�2�^t�=�u��uM&��"�W6�.Y��ڽvu!�%��y˜KY���P�e4� ����&rb�,��u�4ʚ&3�p��r �u���(z��d�R��YW�l��ݾ�Q[��T�"A�N�Rmh7e��R�t@�K�p��͢Ac�mz^���(>zl��]��D�N��a��a���OG���$a�*1�KF�C���M��P'�т�C'J`1�Y�jL�@a2.W�!�G�Ϋ��f�r��YѢ`&鉍�j��:i�zK�-?��q�Ȧ���"��p�G�x�\ݎ�nTcoZ������|r� �<�M^���t�pC�c�<Tvw�K�Lx�S@ ��l`�N����ެ�'�f�q#8I�N��5�gr]i�&[�
JY�?�6y�x$�7�W���ِ_�(ڟ�}��Y�� $��;-�^��p��5���X��}�,��
2/��@���n��~Ì��ت;h�6���Ǟ���k3 >`ѻkc����q7�����P����@{
q"������xb��8�r��F,��K�ï���Y��j�#��(�4bU����Ԫ7}|�y�=d�L��[�6����rI�=,`,�R�sG=8� "�+��P9�ѤV;�|%K�Xt�y#��Q�@B W��F��Ǿ�g�p�]�c�&k�}:��g0��	�o�#��?FdǬ�B���BJ��ҫ��1U�)�[�1Q"����@�mN��&��j�Xl�n������褱<�'8��Su�.8	j*o�Ň��pg����*�+���Tn�q(�������^O�a�LUA��c�����B�9#�Nl[9���O�#�q>䒟���ѤWZv�ȧ;� �����M�L�{&I$���Di�=Y ����b��b!P�c$�>2�P�c�/�s�v��*�,I��9���µc(^?��8�����s�FnY<�)/�/���е�E�8
�(�t@����7�L'�\��xDɽ�~�Î�
�	Ḙ [Ͳ3z۳�'퓓��u�{����>����͖�&p��=|Y��K�j��F��ӥ�78�m;�(��|��G�2����Y�;E�O����d��@���}��qE�f���(�H����2���.9�RWv0���Oj=k;���M?�J���8�m^�Q����ß�}����)�롆x؈�p[.�Zik��Y��:�Ir9*S?B܌r��?9���(S�zi�O2d��9���4��u؊�����Cz��l�\��f����fEA��~��ᒧn��֦�B>�a�rH`+Nͷ\�Ft���q7��!�`Hv
��_�*�.u �*?N������X����}2�?kڪ^��33
(6���[�.k��QNF�]츿Eʒ�~�_�U���ɢ���B��&2��p�8��E���������	r.\�0"��w{�	!��v�T$�wC��MD�_��'	G9�W^��
Z9��'��RBۑ�(�D�4�E/�kMd�&^/��ج/05` �ĖKN�pӇJCnN=f��2BK�nm��8��?M+wu���2�ȴ��M0�*_�Ȗ� �=�'V�߆�G�,��Z뷆�	��K�K��p	^z7������	�ص/=���ՙ�?�`��_��浱,��%'�ռ���8�jʕ�j՝U�N�7̒.�����!�(�F��C@��_�ٿO��;E���A{��֓."~-������)��������ñ�Jm�����K�6�i%���HS`����D�/�2�֭�07�p�Eu65�u�M�j����S������a !��= CTH��f���)��d6�w�]��e$�J�x���Ьt��dF��B}!=_0�%�[��B޷��A2���)��)������v�?S[\��E�7��K�D� �Ek���a�㵴C���p����X䥰��d���7��
��A7�+x_*���C��4lr+廯��YbN�;���(���=���P�<v{�$�@b	+{& ��vs�}��)����s"kn��c�3��ԏ$!3l�'�h�����=3��D��6�;�+kpn5��wĕf��W�VE�I"W ą�_`���a���4��ߥu�K�j�'a�m/K �e�Qϧ�k>�!���P�]ܛ�%|rx�e(�..��P�1A~Y�][$�Oh��m�;�N�7�����5G�sK?�$��D8������{)p��QW>��S N�HN��Z���!����ɋNwƽ��z�~<��-c�$\�>G͗f��&���b��H?�=8�y���O~<�7�[�u��w�5�,a� 9s\N1��������
UGװ���_ⰷ��������$�e~0�nn1&g�pn"�o��` ���0�k��e"Z����X�Z���jfre�z!�@��-�4J6�^����~VƑ>]��Á��za0�ڷ �.�`Iy�zv��=����펒ұ�]K���jJ��w,2�y�3Eh�C�f�;����+�H�͡���C��k��T�Pq�h�1���.n#pݳ�rg���@��&Y^�'� �s���>������v��5�>�-�Cm^01�HjU��s�Ԡ�oM�/I:>^�Ui�舷����Q�D��@��͡in�zN�pBu���K:'��*��x����ruza�a���8��,���{ l]ˏI���po��+6�u����Y����2�ھ2Ϭx��m�dsly+��dYA�R���l+����7�9��nP�R'q!np�N���]��&�����Ӎ��Q����T�3�1#��r��>�<�*�:"+�������d�ISx�^@�'Þ@�ZǍI�0���~�&ҫ�;fsCF ��O6ȀK.X��NوN�r�Z�� �f�c���h���α�b�g9����5�{0��*�c�&(eL��j��%��&��~U��"���*J��fk�^RywZ�#�oZ@�'�����LD!ٶ�Sjj H̇�f�>Q ���1������-_	�Is�U�_B�%m��C�EJ�fX�,O'�[,�$�����O����(�iX���k��2�M����dW�QC9�S3���D�f#*HD�� �{cY�i�����pՔ�F�BJc����	q���c(j�s�\����z�\m�ԄA��� �f�y^�$����u_����ֿ�yN��o�m�G��G#��M����ڨ�'��B߉�v{�?��@�J�ή�&v�,W{��+�R��U�m�jK� �Es�_�̵��p�<�O[\�>�T�kŨ'yz���tȊHў��RZ+	:�f�"Q�0�v�HJF�]{,��cm�=]�6�M�{l]��KA?�^�����6߈��;nn�!DJYOH������4��$�u��]��>\�ݝ�-���Z!��=(j��"�g�Gr�P �̛�YG�F�L�A[;P$��Lr��Xґ���q�#-1��{@���nTn(�k'I��|.Eb�ۉE�f���JfO�v���6d�����u%'P�_1^V����<��q%�WG�*�q�
����7T��q��S몷�}���ȯ0 V���=�6?��e�K]N���H(Ġ�i��	��������=J�5�mk,z�!�D���(Q��ֽ+6TZ�m:����(�1x��LK�)��B}Z�� WW�Ql��\ʥ5�ؖ�i���sܳ8�4+�hJ�$�m����mK��\�����)�6��N�4j��3��`�#�p�&4;jk'�>�! 'U7"�o ��%Ge���H�_��H���8���i��dvr��dD.2dfe`�};|��h̯$���!+��4���,Sy�bR<y�י�(�h�(~W�5҅~rhb�e��Rj���eK�nn�Ju_b���O۔�iL��T¸Ѷ�;~�oD(�a��N��q��D�~-a4�~J��e@�u�1�`�%����';\�Ÿ��2
�����.d`X�%�����uj��qj�@ 5'D\e$֨��[F��K4�X>e�sM9
���{��:����Xo�����,&gh��e%�L,�~��Ď��kj3�{���~�x����f���V����9��,F%��Cv�� 5����E"�C��'�z�ب��y�͓nKb�bjvl��]�_��cXh��[������d�8���i��hT>���<�Z�45C��LӅ��R	�����G��Ko E�Tsk���H�
�`J�-��W��Q�$���%����q���Vn�<In��Cҕ ;��.n��H�x�m������F	&1J	\�' �EI�n������n��� h�Rem`��[��T[�l+� Zgv�@�0��D9J���i���Aބ*T;iGm��?�>O\���1;�c�҆4�׃30�p3�K��`uX�z��n�G����k�H�m�^��9�k�x��7E�:HA��q۱�f��~%|��0�;'�L�ՄBcs'���j$�����W.���F�$�W�ؓ��7�:���_eI��ү���kX� N��Js/�K������ӯ�v�I�
�h�e��9�����*\�<V�Cl��0�a$����W`/|�K��' �G�T���}��F�Y��V�=FK����q��yp��T�>B��X��嗺<�M��i��
�-&����@�tdMG� )�>���2hw����Y"����_u�+��C�O%�Np&l�)��"�q+W��t6�!�>CUՉv^���M�/��/.)��r.q�o^��%��Hy f�g�!����� ԣ�|/��V{������rt�1t2���.ʝ�^t�p�^�V���e�K�2o�]�%�;do�c"D; i������`#�0�F�T��(l;8 ���",S%6�g;�K� ��<�)e"���n�$���}<���D�Q�)�Zq��k�`��~���Ι����C05o0H�̄Q���|��m�R9^ly�#�`?T�|�����]��#	����ǰ���P�dl_L�e����S��H��r�#������!6��]{ʈo��}�}���2�IB�>�SqrF�e�/-eՊ��96���c�}�;�m)�nEC��m[�L�D����ﳹR�6�Z�鯷����3䲘 ߃}[�rK������𩁥�۴���6�cX90n��+�VT�u�n�dr�p�Ƈ�7Ɠ�}�����h��o8HÊdkm�rU:�d��mg�8��'����g��3֨��(jN�D@ �Y�D��Z�ŀ���gy<�Ǡ@�� �|s,�k��@.G��!�6?A�H{hN�įgw�w��8�>��۳���'�� a޸ ���x.E�����ā��on�}f�Dq�b>)��B�{{������
:}�=����h�������j*F)�����-U<��m�����3:�M�2D���n��� }!��r����AN�'�g�l�
�tS��N��~!a��8��4PB槢��P �$�D1��W��M��\�]����{��T0�/����|Z1U�@tw��}��f���\o>D��G���7�h*c�;�/�{�K �����$f/��
V���-�eg�s�L�I�t��eQ�!/먁�O��Q]�ӻ�.���B�������@����(��M9�V>���?U��+m�})�����U��R�}E�+У����vԶ��N ��.�=XH׷YE~��=/��ly1���D=���ٔ���4h�� ��C�%�gkW�<)��Z���d����EJo籡�0�
惜NR)"�X��JQ?���
T<U�b1�=�)��
Вh�9�,]��ϛ驁_N=��m�v�@�'j��٨��E	ĺ��)Q����hV��s5�հ�a���!`���\IC!kHߏk3X��!���P9{1�n=O!w�*7����	M�P������h����Ӱ��g����Y����4�� �r�-��K&=�+P����ݪ����ujs�ٝ	�cMc�q��h�Yw��O�o�Zż�<@0�?����? ���}C�}���Ǽ#ǷiJuz� ��/���?,u����D��i*
��d>��F�Q�&y���I����Tr��Ȇ�N�-iv+��W�oooo�< �UT�Ui�r�3`lEϙ�"��½S*W��A�~f`k7j�����Ow����OZ;	�ڂ��I�r��" o�8�4D�b��5��ٳ�m��%��k�����:�fX!�-@��:������?>�L�_������L��T���l$��7I�����yL7���V���;Y;�����x��,��c}�W��t�	 ؊�uwD�mn�ba�a�ک�o'�|���śV�)y+ ���K-�0��󊀨U-���(��/<N��L^51���L��@�䧾O�ȴ}�w��2;l���0� �Wk*U�=8��)*5���am٘_�y׶җJ��L��xH��� ���n-�E~'���øǓ4P3��?��, 15ե�w�ʳE�n,�:�������%��D�$Xt�V�r�e��F|:,�ⰷ�|��JÏ4)V�9IY�IY�f�1u;�9�,��"X#��.�4oq�2:x��'���6Yo$a��(&�V�>�����GG���yU�G텅ԅhJ����0@�b�5��+N��ɓ�|�~rܳ#Wk���&����5bc�U����;qb�E|a6�[dRݑ� ���s�)7R�\�޾1�e�-����I�T��9a�٢�lᴘ���3�ţ�Vwudl��[���o2�l[������6�/���B����x���\�.,�y5yU��v[��S�$�l�[U��t%�:џ[�l]�,��YJ�P��#�b��8�n5զ �Qv�
�:�d���E�a�/��u더J{oW��Q/���W��k��M���~�΀�+6������	��V�Z
��2l[�BY�z/?'�Ke��C����V݆A�<>��<���+A����;j��*6z���]�`�;�kɾ�{����)f����h���AK���������\;|tC����ʧ�C�bW<�C1�c�E�'����7����钫� ���]gU�L�����
"�O��&>731����y�ap�Shٸ�ݱj�[כ�9���.�ѧc\�����tGr��=[�]/C���Ԍ������a�
쐐�\+��,:ˌQ��
s?��&���L �yq��r�`�UW~_F�������Va�z�ģK:���O�m<�R�J+�[|�x�]��5��� �3��6��3������5S�vT�9s*���:l����G,�����%F-rb0�s��x���5i��6�u/��#Y�ᑍkPf&Xg���b�-&C�Z����M\D
���\$"NFF�}1H�ޑO��w���7�q;D±��iXJ�p9X�"����bP�lIAԇ9��I�^�N
3�a�������c��pq�XV��Y2�h�K!ʨ�F�e�0��ѐ��'#�W���������ݽ�n(!�a����pz:m	�Ǆ���*w��M�9��B�'�����#�?#����Ew��K���39g�0�-�v8b����\�󃺳ļ��n��C-�Xh�<#go¾=��Kyt:Qt���w=��u�j&t4��e�%�+��?wkl�Uad�/꫍��
��G(jX\x�}��
b��F�᠁I����|�'��{�o5H+�8�65���� B)��=�ǀ�����Ǔ"����G���u���O�%����uN�1ʍ����?q;_*=fi���4�?_�*� Q��u��bי %ѝ)}���N����ei�Q�+ ٨�p�FG,�Wz�߃;:cr'��X�V5kvh�5��b�x4�Ke�5C���e����������zq�6D�Jovv��X��������9�8���J�0L�
t&�{�q���g߲�/�������f?ld
��~U��c$!7*�M��v0uF�8������!=o��L �B����*�	�Բ8^����2;d���z�{���b>X/on��GZ�Ӆ�����I�X��G>|>T�rx3b�Tҿ�i������0�{��	�ΣEX73A���_��`�һ�߻�<�S���c����"f\��rL�㍇��͆���yKbl\j��`^C�C��M�������Y))�b��l��(��\�McbƇ�,�k���5 �Wxq$�������8A�%F;8I�������|����3E��F�b"�c�fڕǏ(�K�9�-\��G��K�~��q�D�2���\(�P�]�k<4�� �}�s��G?�z��U��G�=�˗,��S ,��7
-��ڽb*��G�W�37�O����p�|�Ϫ>;ř�ͧ���H���9M�0k�lq2�)�&5������v]:��1.��K�B������4䦠��	bS@ Br�}>��;)}n�r)Fty�4�7�'����������xN��mQ��6�V6�D|C��|K��v�Ƅ:pB�%�{s�E��U��gĮ��Je�*B���g��A���
߄]Ռ���y�HHs"RzJh��B��Χ؏��k�'�����O1�B�ԧ�ڃ+;��GC+i�3c������X�����Rwc�S-�W͍6�+ʿ��q���aQ����:x��;��d���R��)��#���{+���}�h�hf@
oW��Rs���G~�����|��X��GӞ���پI�E��3��=�Qу%rX��♩t�8�.d�q���� ��'%ۙ������P~���̮�<�^��>n2��#��	<����j���@]���y3�Bv�X�N����Tɡ�bJ���$�iXkb���S���Aeu� 9B@!#��c�SɊE�z9�]Q���S�U޿�s�CkD��Eq�uҒ�쁐ls.s����K�~�m��nQH��u��C.M����/�@� ���9�٢!}�d)�_(jɛO�Go¸8?� �C�E�e��0����R��v�U����l�{��Ļ͒a0��Yz�qK�׺�Cwܦx���F�d� �>s�+�Хa\	�7F���h��#��A�,�^6z3����gf!|4��A��΢��
��T�j{��N���n��{��٤��h$�:9Cش�8_�m�v�ᙙ@�9鏡�k}��XЎ?���X���OwG2>:7�:<�o�����'��V��'.p�����aU���B*rl��:�[F��M��c{�$J�m��iS�a&���\.����u�%��"3O�@����t��.�j�k���o�H��?ng_ T|x7�_�(WN�tOJ����v��J~�ص�[n���;F�[w�����cJ6"�xuK��i9}H��^n}��-��MI�a�-�!��ka�Z��*�vA�3"{>gjV��kȭ�귉�}i���r2�zFģ�)������4�W�9$�T𹒋H��%�(
���Q8�D88t�e5���dj*F�r�yg5$������(�P�O0@����r=����aG�p'j9ڎC�wWq�= �`��#� c�txZ�hu�\v��p���4p�7?%���I	�t��[޽�x��R]�L�{�����Ԁ*���wZrn �z#Y�i�|�>@lq8�QC�f�/�6��%\}�׮�M�|���x	���빱�x��g`�L ��e::@fm��'��w���s��폜��I�Fށ淮������[	�y�s=����p��0A4!S+�c�>��RV�]�\Y-��6Y^���.�e�|���^�)�$��.CZ�<�wN
�E�e�:�SRH��7��=O�7v ��J�� ��W�������́)P��H ���+��q*�P�Fwq�������,�[pɖV�fp� ��`A�a�fJv���L�@�V*��E:9�e�3��Y[G����ż�� ��%��`���1Z�f��������3��]�[}�7����"*�:�ì��(�]�\�\��>v2�·;u�5�K�o �2�F�SIR@!�z��Fp�G�@^4^������2�O��q���nn�V^d�aSX|P���%Q������%�}��ǉ����a��H�\,,"|�����Jx4'UBo�*w6<2ɳ+�+~�q� �Ϊ�C[e9M�A�Qi�ϭ+dpsk��Ȏ[:M�B�f~�{	�tW��=��ֳ�{ ttR���
��2����<�!��,�2�#����M����7������ٝ�j��s��k��S��#���u	C̃Cz�W��>�mh�1j��ǃ�\�n�tN1�6��}�c�)��l�{��0Q��38w�I |�v5&�ں�+��T�Jzݐ�	��~wE�����o��Y�Wm��p��{��������>",��$���{.]>�rF�I���瑖%���z{�f{=�ņ��G E6�}޹���π� ��[����P���h�җ�ￌ��h7�Rw�����z����.�u�'�����%RN+]*�ow&3fϸ&'��S9�k��UVs,���ܥ��`/�Y���t�{�����Q(QU�ƕ��+�
t�F�eh	�v���Ӗ�U��)���@���ˈ�f�Yχ�E,��˄\�*ӄ�Y���/�@