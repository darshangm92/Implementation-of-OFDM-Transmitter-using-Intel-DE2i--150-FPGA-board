��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����胸i�J�y-�(��*�U1�OA�7�-��/��it�Y�Mv�}˽�L�:�^G�U��/�y�
�[fz������ �G A9�+҆���
�-����2$�6>�#�̼wC���W�^���D�|{����˷�0��KɠnBf2�3Yc���6��T*ɹ�~菚�JsE�B}�������-Cs%�} �Þ���7���f�f�)4���m��֯�oR���"�;���4e
��k+���!�r�S�Z���¿6p��]j���V9�+����<�I�u�(�C��7#O��_{����ᖓ��n���8�����*�ho�	�E��;`/�4|��ع���`���s9�~��h~ �*N&vo=΋��R����t<y���
�dL{Ȗ<�v���I:�`K��U�e�<���T|����C�im���CI۷H��%⋎����f�(iߛ�� u�]';S�mJ�b��k)�@�b����V���j̆|k��'�f߬�iN%zcU��p��z
ɬj�P�yhA�¥�J+�i���v��o<dՌ�ϖ'6ubט�`v$����-���^AJ����S{���NA��� -o�d����s�O��/8R�f��s��h�&�+8��)��:�$[)��黝�)�u����M�1�S��j~9�s\+�K�������׹��5�S/�朘�o�tI���hCyȾ+�B�Ō6��0�?���o0�"���1�T�����b1A>�a�_z市I�#Y @��xDV�� ��:�O��~y�o�#�G�k��ah�����,��g'�p��X�ѥK����vx>>��伳�^�����;�;9	�E�'��'��$76\��1��ϑA#�	��?2�3Po��?�0�(��Y�4z�؈�����w�����G��2H0B/B"%����)�LX�oX��z�״f�y�YU(L@π��9iD����[�RN��<��
έB7��_F%�|��:�����d�$�eJ*")	I8�����:3�T��n�,���gA��؍laR�%��⭥k�e�#���t^��C`z�-�����M,�8�r�܅��I������G&+���b�����Y��
@ǅj�t[)�KO�H P�ޜD9�U��[���Z-DA>��L��"�e�G�T�|�SL��m^�k��KZ�vD�V��z<4�'�w���h:�%��;�՞R�����3>D�@zA��挄V$/��^�ո��^�E���C�N�'vr9\�G��l�ɠŖ���L�iv6�_߅#-{�1��Jhҩ�?��'���[��/����V�V T�]���f.ˉ���<`Edx��ѼԭY���0���57���3J/�C~j�এ�8.EQ�V9�y����T�IC�eoh3[���ګ�;A��=��nP�1,�}*���N���6W��="��B�+?ֲI!Ln����J�M鵙�k�h/s�-�Ɛz�?%�O������|@������o�N��ņ������J�� ��> ܞը��5y9x�w̐���F���m]o�L2���+���vLU�Q�4���cr؍���7qW��'�8J)���J�B�Z�r0�76��Γ��U�����D���%�Tu�^�b�έYq�E�z z'2^����O�.��yē	Zgܥ�)	"<jÆ��Mc��u聢���>�׉F
T��O ��ڄh����
�����<��#�*8Z��w,�Ol-��V�s�(>*Z_��Dky�T��w��,L���|G)��{���B\z��$j(���֯r���¶�3d%7�!�=mk-�|[��z@m�����,�;e{�mit�����.f�
�۷�
4��
�;��-�֑�M��W�.v�}��d<i__:*rkܓ��0�F5eLCw�L��{�BW��4���v������ll�o�>�|[L��sz�Cm��������2>�;g:$jW�=�Nr ��������7|o7�4̔�g�r=��rlM��Ui��Y������`C��`�@�f��@�{�I.
j��NȃyS�a�&�Y�4(G��Ǆ�!�.��[SF# LB���*�:���������֍{�d���,�C��+Mq��D�Lg��i�-��Q��{W�U�f~��Z�R)�P{�P�'�ٸ/yN�fFS�#�T�C'Yn��2n�oh�u*�[�`L����}��?^���xi=;Rk^��%�<�Ss����R�NX�6�I/�!��\�n� =�zo�d�K�����nhT��M�_�����3�=�dA������i^`2�G�}� g�o�&+�(jsP::B�z%$�u�ׄ)2��^#C� �GTwb2��~H�UH����MZ|�k�lͣ���˼I{��Ǐ��`��}�9�L�t���%�p+T���9|8h��y�q'�B���a�F	��g+Mnr������=�F~=��G,\�5�`f�ki�*ʹ-&M�\)�{7�$Й�_-�G*���ŋ�m#����_I8��CW�1n�j�ܐ0��Tk|��G����]�0�#U�!�D_6F�����*�k*�[�
��.��,±a�Ř��^k�1rU�n��߲��6&_y���}��ꑐR���1������۟\�%��D�V�F��� ��\kב����Uݸ�� QAз���6�$H�oWOg���:�*)�Rc��a%�	\P�o�{���q!Q�{�pʧBl�=�Pv�r��d�Oz!�@���M��[-OXq�ki�$@�_J`����~�1BI����C�AWlH�I9��π��x�>����-�҄��� ����O��1n�l������Q�����|WZ Cj%&�o^�5�b�}�m���؜7	'H2;�UI��i�����|���:�`
&�L�����:'��4� �t6�j��[�:���[]���W�"��'l����sz�ud����^��-�Z�����`mK�1�,�6�������@t\#|ְ��6�vg�"u�
���0��㪨�kAt���H��
�7�8`<1�Q'q4�I@�	�Np.��?������Ҁ�6���7�����u.2�t8r��4�I<(�'����?ǰ����L����-�6�w
7��*j��>qo��zֺ�qO�)sct�h��\j2��F^}#�0�a��(�b��(g� Ņ�w[��2����zmML|��Z���(S���,Z:>|��c�l�&a����W
`fW�08�)�L,3�*�����fo\�
? �;ː),ҲZ��Q�2��c��	�u����r�}$�
�������Y��?L��@�x��������N;u/���R¢��qy�}9P�Sa[�kw�uH\��2��oɑ��Ӧf3�2z�	�{�"�U_K��w�`��<��3���}9oA��H�}��"�_����;_�eլM�!�;4��t�ڄ�"E�1z�V�)��X:?�<It�xZz�
��K�WџZ $�����Յ�2Z��b���#�i�3�