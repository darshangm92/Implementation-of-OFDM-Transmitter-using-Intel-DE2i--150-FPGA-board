��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����蒋q��x2��+���Y=�$�FxV�q݁9e�^v���U����~�����:�GG�BIF�,�r�a�BW����7�Z��z�A7Է#_L���E��a7 I�hn��.�!m
J��[���~���.�c����Y��	g��.�J�
l=O`��p�̉���	8L�=���!I8�f���)�&Ya;Iݳ�UY���}c i�З	j�"�S���F�踢��&K�!����~C:%3w��� �A��7j��h��S�za|�3Xv��k�g��;�T	J�+���L��fڠ	4�H~mq%�$g�9��K��T��*��PǺ����-	�$���Й;s�0����F����-ESo�"\הXaP�?Ѩ��7r5G���f�H�<���a��-��Ou� �u�đ���f�'#M-{Ѫ�8]X��n�7Mm�^��)�T���~Vfs+�r��<6_`ƆW��t,�Uظ�+M���W��*��qخw�4Cʡ����˿e�o@��Fr/{b�[�l��$�3�\�U9��)��
���	#-MJtw�<U,�����Y1C�k~`�0XF�a'>�슗�,��aS*#��Gx�X4���M�W�O�����kU�(���g���j��u�,�����0׋k�A�-D�U�17;��I�.�d�E�h|a�1aͫcfԼ���A��p�nw�����CÈ���s��D��zr�]gq�_���1��!%�"Z��%R��a�}�1LSc��9��B��.}��]I������������b��!��sOp�U��$�AvD�Q���9h,���V���Ln����B}8�F���_W�Oi�2O���o���$�hom:�BI�)_d�c�K��������k��͠���4|cD?T�*�^_I��r���1��Fˋ�i|b `#ۂ���&R��'g�<�ލ��c%#�;!'F
�\9^��<�=�V:'v.h�����5
�K���|lR"��xf(<��.�QV�=��E���}]�\'��Q-�J\�� 	T���Ԃ�T3��t_�ҵ��^����g]�E�Ͽi�j?�st�텿��4j��}�˧0�,�p�ro���_+���bR�Y�d���<rd�,?�|e��2:E�؜ٴ�i�/t���Q+LϠR���5$2���j�},�"g'ul~^��W(�,^������ꁆ�Ś�e<N�9�hv�>��Ny�a�����>I�	1�%A�x�gg	�ǘs�n����~Z��%)z�0n>Ĉ�.��	������E�������iM����7�����K$;��M'g����\v�VkLF^G�|��.,4c��1�Y}r@�i`���ݺG� |t����롰���:���#��}�`3�T�&e�^(wG�$�lWU�?���i�A�I\G���7�[���9p�"��l�!�|3��p��eO*;+���Mn�V����D˭cL����il�&�P�o*����8;���N�D9��52��1��Z���DzQX��S��[�Lø��G�E�7oΩ�A�E�wEg�v3p�`��J��X��vJ�&-D�"�\z��
�$Ķ���"6�u��p�<4,���o�]�|��U�=�wm�p���5�p�N�g0Qsث!&�G"�}���(�I7��b��*	e�����L�t�aK%�h�S��C����mc�}0)�)�/�+6��b�|M}b����}����������t1���RQu�ދ����,�G�Yj�A���>�S��Mg��R��ٸ��p���ľk���*E<��U��"O<��_^��4�ݧ�@Cx���9�@f��xF1�.�^� �u��c���������ħ�Y�XV��zocg�*���|O8�r�/�������c���}��L!��BwNOaR�2je��]�^e*�Є!{���횧�����fmMy۠���a���;�4����]?�`zQ����i���X�0�Q}:W��B˒sx�DgvY�����T������L20	sfЭ��7_�g��C"�����]Y�4q8[�O~��wM���C9ӕ���*�G�^� ��;������1� �r�7�\@��S+�_�b�s��8�su�B�TYl��Z���=�	�ΫəW/��;q�D�3+��Q�����lt�~B?��k�P��B�E޿'-CY���d`��[G��	�������w���i�E6�sg�� �����^Ł�?�q�����d+3�s��r��
�I��n�YM~Κt�Ĕ���ض�R�+E��m>,b�F��S���TN�Cq�����f$K��K|�W�C���U�Z�4��~����J6�U�f��F�ɬQ�N�%�#�晴����*��o&��"���.R
-���g���'���*.yy��bZ\$*7
�m��ѐ��(N�0�'5��)��Tڰ���m+��x�����o�� G�ad_���
��Q��gB�Ӻ3�91x>�io�9�}B�g�F��:����HdAt��9�HG���BԹ�G���C͉�m9㾈[����DT�Y�I��`My^R�:���}�.q	`C�&B%C���O��7���ҳ��:�R�C�6�י�'M`e�7&�_Q|�h�m�ʏ`7=�z�:8#wO�nm��D�c�0�n��r�i�'#���6�H���W�t4!<O���]!s���x(��'��	�4Q��xBZ{��&�2��0��3���d��<&)���2�`�z��4ڇ_����[���<a?���䳫��%i���C�HE���p�CU�|��k� �}��*+xj�Fy����������I��9����J>-��J
,v[S��De�IC�{��/Ӗ0;cj%�,X��x�N2�k2�x�Y����=6��"�W\�^~��|a4gh	18�{DJu�쐂K��ʣ^�����Ld��VKq
�M#Aw��r�#�k� �DSX M�
��Sz���i�'w��ՙ�q�͆v�n}�YfKn�}Ӭ�䮷�����$f�A�_"�ҧ����>����W2#��w8���9�	�Zae��oZ��5E��:K4zmI��oPw�VLon4��ŌW��dT�J̝Zu�lݞ3<U���7�RlH�KX�.��I2W'q&"涱�*.�к����h����c�t~����ņ��v����p����3�Wm���s��)�N�A���v�K�q�
�"��~y|��Վ�$v`�7�6�4�7�CO.}��(�#ā��5�E��Lӱ?�ഹ�e�<��T]G��w� mjE�0�4ӄ3�5�9����y��5�:�I~� x����} ��o�v� �+�:�ys���k`����� Xv��/;�TW��S�P�z���=Tq �>���8I��Q�ⷝ��2�y�<����9�oB��1�ekI���G�6����u:��"�ņ�<u����νW��n Vsf*65	�Βy��T�ky>��H9�0�4cL�Ϩ?�1����ΕI�Q,�eS�!><&�Ȯ�"�6>���o��s�h'�t'���k��o@^�	�C�Gn�喤���� Y�^�OϮ)&a�+|sc���>�K��t��wï}��S�|��U��d��.al���pw���CA���t�e��~�҃���(%k/O>nz��Vj��3��j�/�,mZ=yt);+.T�s�@��t��y���3L�?͙w���,� ��36�v�j�4�\
��v5}]cD��'�5C��2��sϰ5w5��s�+�;B������,Lc��+��N}�P��F@�}Ψwm�g�GJ����I�ny�F������� b� ��D,��h�^��'���m�����i�y��8�����*���*�t�H5�P2j�i�*�u�������	�xS�
j��m�	�?	4B�@Ю� �}�Q���+0�c�N��LM�򗲩���Ȧu���K�e�>f��Ǐ��#�
��t\^�G)>��nB7OՉ�/�/�s����5q��'ZQ͌�:t6֢2����E���I��(��k8w�+�����d��8[��i����ܶ��"�F���xl�{�k�J���/��f �"YVn21NS6,�Q�3��ۗ�)ص��X��o�K�d�Ǵ��mi���������������k~)4�ᕴΕ�_9�9._�h�Dj��uc��B������wٟ��D P���/�ځ���L'k����gs�`�·��nrm9�5�����2�e��Y�� i�fT�%���!�u2�ب��k�B@�M6z����yB���<��_�ȝ�vhn�Ԙ���r�i�>$�L����s�zET?PP!&�OXk����|7��q����\h�����Ԁ1��i�C``c�l�R���C������@�vVx-_�m54[,���[�ZL��WJ'0N_TE<X��2�5�"5,�P�>�;�;Th�k�|FP��.��$�����R1��C���<�f9��5W\q裬�q��L���~�1�f#��@Ж8�/A�0�$�)"op�NB��L��^�yA$������k�S+��v��rBٽ_���}���4��a��˧���E ���h���� D���cy���vM�n� ���y���b�A��ު�[}t��}������e�{�����]p:�ߒ��lr��`�ML������)�}\��a��ΰ�;�X��`�@a
eE�"(fuT2j��/_��Ԡ��e=�t"a�+��}��7 �d�t�]��ր)�x٬l,�ltx�7i�Bq��v�+��i�3�H�`{M;a�dL��SpD|�vu�eI�*vJH����G��5�B3��@EUD��i�p�<)o��}E$#�;
mj�j�,Q�S��Q�)��{}1�����6��Ы�5�h. �C�:�r���BTo=2�v�Ll�j-ӈ��c_��t�������a�1��c�/���n�|W��Vᝡt�T��:}Ed���[��JxJ|�Q��#�=:=^�nRܜ�s`݉T���A~8;݊���Ҵ�f��y�n!���p���
_�����a�RC�>���'ٜl��DA`!k���h.��S��VW���-���u�+�)|�̰��G��\K���g�aU�����24%�VO�D}:z�������Z,���C_0��i���%Ic�6�տ�-C������:/r]I���7�]�˽��������=M������[���F��� ˂*i[�M�|���F�t iw�m���2 o7�D�&sW�t��>�#� f�i��ԗo�'���m	|�s\�뚐�269��� z4<s}�OjuG$F���H�#L9�"�z����sE��S��>��~vC j�5���<����r� /Y���\�1�J�E���'�������"�&�gEj}�a�V^�����'�~��P?�ۯ��X�"N #|->��p�w��x�r��a��Ux��'�Qu�Kd6W	����;�E��ٺ*�֡_�J��H��ܒ]���=ȀYP8 ����A}�kB�'�x�H����	By(��u>�<Ï���褀MV�X���:���M}
���������zv|���
��}F�ܿ=?~)k֘��5�ɰ;a��d{����!p�+��f(Q.f�P����G��թ9[B�NO--��HK�(0�0�,�v�xǀ�%J��PI��?�3 œ3����"ⷚd)���#e��{��QW��d cs�h3��R#����e*��aT��	o.���*�i�ۯ@AGWX����=��O�p�TZ��r��^�&�%?��0{Υ�x�\��!�3�H�˄�q��8�Ng��#]tܘY�T�� {VnCC$�K>�_6ڜs�y�$$$B@TP��)D'$����SS�Ő
��XM��T���J��j&n	$�#m�&�O�Ę.4�)SAA���D�Gͻ`Kǂ��g�B@�6��|�2��4�D_�&]�|��*��5�7�Ib�SM�e�C#�Knag��� =���P�#�B1����J�����!�7�Jv, ? �-���ȘrF�Y�����彆�K�q �� ���N�@��e�1M��a<�	1�z���R:J���	��_js�x��V�ar��k���w�aǘ)
`m�1��=���~�����$є��G�w�rT¿4�0bb_�i�gŷ��sT"�����%����^�f���R؊D�>R�P��}*�$�,�X�Z�pN9��ѻY��o��1�z�U���zZ�2�e���|n?G:2�(�K��b��}$��8|���DJ۱eO�R��S�4 {�А�͒���U�[��	�l��Z�U�%��&ť�'R5��O[�"���!Jǳ4��ĝ< �9_��*ץ�+
í4�x2F��^S��`��}�������pF�Y-�=yhܒt��H)�J���_f�r2�ϟ1��%kJG"����m؀S�kteBϸ�)�r�C�2r��	�p���v2���aw݈�8*�F�j�����W������1�$vA�fh�E�B���c��I�ǘ�B�ȸf�������yv�&(s;O�k1���@��^C�a���N���"�ً��1��U���:��XDs�kOdL���T����('���.�\2�Z��U�]ʉ����M�6��J�(O�q��ʗkg��jIԵ|�N:�u%�������1�B��Kk
��9�r�(�ժ�-�OJ���T�H��氧���D�ª�y�}�8H�C��
<��4 �ߒ��Z�[/܄�[���)��Ҧ,
�+��R��O�_�v���d�~'�i�Q4�E�1|�r�NG0Z|y������|e��]�E1��#50q����h�AKe���֙��
�=���t���y%�2lu�������M~��k�ڱP���e<=j5�>�	��9
�6U��cꂰ�9��S˘���T��6�{�0c͟B���<S�q���9��8y& �D��|Cᗎgw;ٮj��"7C����w���Q{E�͒g\њ/\�j���G�4K
��ُ������<Q�WD����1�5��Soo�bS�!u�rp-��q�6�����P˕����s�u�uQ�^0c��x'��E�b����2��	Rk
w)�"�r��d9^e6 �=
��%��h!��&��a�����p� ��kQdO[
�4C��	�V�Q�����J��I�҆%�ӟ�3��P�2�n�vDI��%%�����i2й��O <~�[��$T�{Vo��J���"Olkжr�q ��� Łh�ł��L��jJi��C�� /�q���[�#�<R��.��/F>U	$�3?��	�ǋ3@�z��-9�L2�!W�8$�xj�D�����XKB֫��D��d�[;���Rz��X>ó���k�����sٞ��C�?MTi*�$��i}ux�3p������+���]��yh�
�y`#`0N �7����S�m��O��p�Y�o�L�w(.�4@,:N�1�n�[}���DF��]-�ѫ�/i�K,P���[�f�ar�z����T�-L�Gcg����d��:k��gM����3u��BXϔ
�;��fv��
����H`l:��0:��R��B�-}��_��/����h� #{r�=yt����tĢ$+~.Z�� ��&����ue�Jb7�'�2�/��2� 딊��G
�A�Q4RG�|J���?��t��Էy�h���f�
�n[�B��2��b
�)�b�+�&r�:Sr���0ΩW�o�3�b��Z&x��R���:���Vݯr+⾭~!d�gu������Y�P���I��P?�ܯ�hV���?�
�c��g� ���4^5���]�������kdA�y��w����y��Z�9�����`����C~��"�J,U�(�Ţ��e*x���c4����#_�6�z�mR,W��i��hM���G�8h��������I�����Gm5&S
����^qT�ʡ�]x��"$��¶�U6��n��P$^o���KA�����:�_�3P�'�殽}�J���n>����"�}%1��c"��{�_.����B4N����ǅ�=HTO��NI�/�E����5ʘ�B34�g�"�=�f�JVD�|_a�6��K��*�7��6�o�Q�/�,�w���TΨ�P*���	6 ���Kw*~�v���܋��U�ƶ 2�U��u\��eo2y���c�}Ƿk
߂�,���?i�ǆϹ� � �ob����/�!}��
��_1G���h
�����t��>�e�"��_/e�
0\�UvK�y��m�����^�į�j��1kI��9���sZ��PJ�6"�������+:����!�iK�L��r~���#h�e��\�PT>�$(|��L�����R����[F{H�NB��S�z���E:Dw�Ԕ��uD�9��%�1�CU����@��iּ�[v�h�AA�}��Dw|-%s:��P�hT�%4m��72&�zH��&�7U��\��!�����N/�bNZ���en�	���������oaK*�SqD�/����^�/d�/��Lg:W<�pL9o3�@l�`8��3iCNQ����Ҥ�	��G�2&���v��JGl��M:˲��3c
�ð#;
�f���?z��}? g��u�	{&�B�<��T�� � L2 �ig�DhP�k��4�D�N�]��3����yTG�@l������Z�)ù��Km�gh��,W�Ê�#�
3lo�B�O���9 S���:��U�Ia�{�6'�����	�����韰TqvY���<ui2�I��
auZ���\�Ҫ���ˮk�rz&^�@�4H�|rS�'���s�-0�{�a�$7#�K�֖��&��4�y��%����=�u	PRq�Ĥ�1w�ّڛ�o�F�����<^�����RxsYj��tOI+��&�㔆����җH�!����p@l�$C!����]������0���s0e�k���ޑlδ�A���P�����BX=h�t�;�����R3ĩv���"e���C��+Aٱ	G+cc>Zf��J$��!��yڛ,�������-��Ҟ���$:6	���4�)�S�w�S�3�f�8e�a�4��,�j_�Od�k�iT�*��皲=�~��S
�vvD���Q��7gQ�u�R��S���VlHp��p��q����GN�]?�KܳT�e�� �!JzV���Fcղ2�����%��%U=��P�"��K|�[���[�����O6ucڙ' ;K���_@3�1k��q.q����*����Y��//�VP�Aaj0�nN��A��Z)",;-�W�bu�;�$�V�y�I����� ����b��/}L��ts?t-�<|�����Rf�5,+|)`�B�Gڒd1��Iqṯ���Cvj�K��O������[�O�5'q+l(�"��Z�����
kk�l�t!<��*L�	�|�?�H�#
�.���Y����0��%q�����.�5������6 ޱ�;f��Ű�D�R������ٗ�Ue�a��p䄉��Ea�N}�?���I&9xy�ħ˥C���!�CNO�LL2rȒګ��q�����?���귍D�A�=����^������o{)��Kzr"�A/ȫY,a#�E����^��7^�32����ntEr]q�%(ia�_i=*Ā��D���#6)JO&Fw*�jr�/�3��6��7Ӊ����kTǵ����י �}��ʾ���0�,��N�Oϩ��2Њle�,��$��A���~L�M�
���������뭐�������D�鿮��#$I��AXѫ����$\Db\�5%PKw���{���u/�mјMՎo�Y�	v�Ϟ����Ƶ�6|�5���aB�i��yۚ�[soG�/bu�ˮ�d��|�k����=��$�=��{0GWg����|�8����J��U�Kh+������7�ʁ�s�OG��1�BN�r��opt���wkB�����_�q8J��w���v#���u��hT1~߻N�s>�>w�����
 5�o�?�4+^�ϰt�Qs�!v�`�CX�9�Rx�?����|�\��HW2Y���;�nw�?;�u��/��S6�f&�.*�qO�8��L3r�а.CD�ƭ�K�ILV������Z}�w���� �%�O�r�r��#��ȗ��X��XX�_w��u��Xw-���r*�{ k�	K�E�6�c��,{Of5�{��a/��ە�wC%��
g�8��`)�Ď#?½p��C��;���,mS�s!��s�Z���W<?�Bǃ1��Z�ݴ������f59~�%g�73%���X`����ˡ�	�S
;��[o��Z����;��gW-#☠�<��N�J��R�|�$7p��sJ�l�I<[�~�>�z� �Ls��5DP�ѻ�=���ŝ�kW KȝnT�Ǭ�o�����3��ܥaR��j�=�mi��WR�X�?�W�CI)V�v������_N�e��Y��Y�A��"� \���.�5!V �M�']����"��UG&�$x#& :v�<TJR�n})�l�Yu�
�Xt؝��o��Ȉy��ҧٵ�����>up�ͱr�j�tʩlAX�*�)Q�1�!��pR.�U�O�g+;|��Z�D�?��-��w]�Ci��鮽ťa���A����ϣ,��R���>n�s��GZ��[��Y���oH#�f�^�L���(v�6��m�(��R�6�蔗����U�iI
��fz�ȏy�º �&jpK�D�#g7����e�c
�������x�=��ũ`�j_ݒ(R�\�Y��k�{���yU�%M��z
��$Och-	��n=7�qHӁnn���2��)�U�wG+r�D��/����L���[oa7��$�Ff�[����R���r�Y����χMQ$�c��Z��,�?���tI�OtR��w�q��co�<*1���jK9q�W#�+�xQ�]y���
�Z�!\BK�S������B^��0BQEe͏b�ʛ�mcl�#������I��T��7�+P2�9��w��	
Q�\9��{�E�v��T��ǅ�KF�iɀ��_�H��O�\��m	�l� �Ӌ锍�d���ʺ���m9TU�%7o({� !�d��)�X�.wKT�!	J �wfD�7Q;%bV�-�e��~�?��q��!��F�8�X��*qĹ-7��[t�O�'�˲�_pHf�"�� 6�De^5�--f��5@,�*�$4=�,�����E��	��A����Qk��D,{`k�nKc� ����XI�&����6���kF�c i���|�9�� Nh���1>y%%�F	 �b3��E4�=W
iP��w�K�����O�_ʰ���;�^b_�`NT3�WDïNE^]�a h����W��$��U�Ɯ�`��D��Kj�A�`��
�͗��im-�b܋���C����|'m���4 U71&�.�zs�m�~��>�&T�&�����]a��az_��R��0#74ڋ�ʛ��1��� ���\�Ӯ	�JL"f�sB},��/,�@b-+�!)�G�;�<���q}\�qy�7:l�V���G��U�j����b���h�4f��hUEY��1!�H��E:
3�{��m�hG6��wE�{Dt&qHS�APs�t�8.����E���T���;)
���Ĕ��)t�@\҇AߠQvI8N'@Yy@�T���MY`��ߵ��m��`�㋆�xK�ވ�u�#����&OY��/���j����boFS����{#{	�t�5�h�s.� �Vl��f���(R���c���o��q�<����JI��3��_��P��%��T��j�����%,oa����+�"���.G����Z��H$�Υ\�#������ڇb	�cB �V��l(����NqB�/��m�������K���h������k��x���;��
��ph��+:�bX��{��R��:�Z�����ÚAS*��əo����Z"�!Uh���T���
���������?��� ��E|2I��Tr��I4n�]�E�Y�؂v�ۛ��/y�e^5�}���&��C6��|�:'C����.B��ǜ� f�3�N����n@I����O%5G�x<K"�6�>��R�^����� f�8���d�J��*��9V����9O��N1S� �x6A����V,3�7�~��Q|�L��{��TBM�����S�ʰ�e?}�x{V�@=�}����Q�ϛ,F���G?򻢸�*pz�%�D����w����^9Wq��<�'�.=@��݉�\���Eϝ��=�oY��-Y�4'`jW
��0zs��226G���<Q�ϼ2�������.f6�p�H[�����3"q_;Y��RJ�5�t�V����J���J�)=��u/g�n$U�TͶPc p:3T �������'+��Ԝ	.�|���Q�G!�J$�v9�M�>@WP�T�@#T-�9j�JI����H7�*�sL���AWČӱs9"��L&,##-��})�Č�*oZ�W�[gR�6�c`S4�u������ʻL�r�}���|��Y�?�w����be�|���]��;_ԐL~��j�r�%ޖ�p/��2�g�����W'W9\"�y3�����E���Ը��p����;e��VRۚ�����������$��˃�f��Ň\E5��h�~�4�#'4oz�4�::���(? ��@`�x�tז���!�IZ�+���M�!�[��~WY�},�a���H�C����>U$s��l:��H�����Im1�M�GWbl�I����(�=�����=��Y��r؂ڔ(�e���Z�K�;e����!�F9��Ұ����so@�H��pJ�����1������kmU�r(td�6y���Y>���RI���F$i��o�ⶇM�5�jn�/�#�T��� ��c�(CwC�ls�\a�M�AJd��Wk<�a�1ɴv������e|��Zos't����Q�����M��2&%� ���+p���Dƅj�d�)���A�hsTpwca��D�ĩ��ֿ>���PV��~�[� �(��?���Og�!�0-�XK��t��R��K�1�N���#c�(��*X��5���i{ vQ5�{�ַ�I��u��G3ET�>X�	"7?�+�μK�I�љ���/�M�t�y�h����?�'#s�h���A:.|2b��:0�5)�_�
�P�/��u�����7�&?�{�	�_o�\�z6�4�5������)9.��z�d�;̢�d0A��3M�[Ȣ�E5;4����O�qR���!4pV��mEr������Ϋw�����wkC�%{�*\Ix�Ѱ�w�C�[�F-���+OՎs2G�`�?Zn��=F5D�:�1���|;�:F��Ir��_���3��{�)������W��
���K��,�Bo���[��ɦG6c�)*��݆�}�����y����{fh5��ב��TY��Ϝ[��1�r��Z#$8����P�=B3]�4@�̎���@������)Z�.MR���.�jF�YE�T��ש�f�t2`b�����l���SLA�u`NvM���A�����=	(	��|4FW䠠�A*��{�N.����܋���_�L@3qk��'6�V�x{����R�z�#���>}DB/�Yx���P��S+'���uFR:��2�{�1�V"��;�!�H���ҔP�'�¿�=�n�K.�;��á�`K2(+���n@@u��H���7��L4�7��N��>�����G��ί�^�V���x�_%�ʰJ7R[~v�Ӷx�f���a�$�牖�.�W�v,3�}ί����S>C�wnNzCx���F>qHt��������P/�-=��\�ɞ	a���H!�M�l���I���6��+1;քvz�y5� u�.;B��X��	E��?A�2 6���.��2���7�+|�1��1�h�l��̙E>�#���f�F}6��ЛA<V���^R&^��k���ohC����=��М�).�b�=ϔ�KN7��eP@YS˧�h�#��m�ost:!T��;�n�­� �O�6�Șs���R�q%�0��h	,m��ъ�/Y����Y�a˃�֐L5�j���?Nh�OE�)	�\�=�¹��63��\�&(4,���r�	)}���F9�;%G�NK�Vz�h���b0n��b�)Q�Ft�[�e�������^s����7اY{�$'T(�~YTU�5����fc�J����"��;趼7�0O� ���
��?��9�����z]f���y\���u��˱�H'<�vG��~Y��- 9K��,�փB\T�tx��)�i�\k)�J����3�8� �9�t����9���D
���Z� ������y՞� �����0 �_��}����psU����f�x�bQ\ ���H&A�Z���z�����Fi:��e��욱e�0V��C~?�X�G&��cu�b��6t��/�j�Γ�ŅB�I����Q�=��9�/�9Rh2y����S� T���I�]��zb^^�@��CD4��k�%�k�ժ4�|����ޚ*��q��
��r��ƛ�$�߰AS�N�O�S!�����r.����E&#�`�?L�;�=`�ZW��Մ�N����(�,���[�b�����Ef�ӏ�T&!��'5c�%X\.v��}f�p�6|*���=-��<��Ǒ�����=hH�n�K���A�L����y|`S?,���l<�w��I=�U�X�RY3���OѪ\�T,�*R$�p���3TcJ[߶ܝ�?�u�z����7�p���o��,k��b�7�3�g܆� (6����"z
x`����.;j� ���Lŵ+�~t����̀�kg/]Ӥ��_w�0�)�%Ǘ�O3&����m�B��Ô#�����U2{OO����:ժ��&��a����8��l���#*t\��ж�}���,�>t{��J�ݰ�ֲokșU��<�ʄuǶ3��v�����>��E��bk��E��X��x|X�}�蚭	�	d�h5����:9v+ih]�9.�Cؕ�E����\@�w���]\������2�WY��)�"H�@'��n9S�)P�_	kn�whؙ��V:�_��FUT8�3��˸qrT7�W�nh��-7����r�|�c��̭n��E�S�r���w�4ث l��Jt�n#�t즆�+2
Q; hM��k� �y.�`�O�לd�4=�#��Ќ�}BQ�@%�q�h/0=���X��������<�G�X��bR�^���~�6*W$��K<��!ڼ�_-8�2��i��!���ݛ��K~�@���H@�����W)� ��_��nzW�<s����J�N�@2%k"`m��)���л�Mu�xe��$A}�")2Q_F[�� ��LMT�ZDi�������Þ
\�OY�FRm�cT	v5Vފ��2�Ն����k�n>ӭ Ee�m�(��_p&)�WU����� !
(5��~%�5��=�7�[��=]��%'z�=7��]� 8������QLVC��['3��A�i�=����`Q�$��ޜ ����]�{����R+���kA���<W��o)=�Ec�FS���<y���>�;���f�G�,Mq&o����4'*��$����w1�	߅jõω���(��5XCIؼ?�Ԯf��w*d��`�P�W����{���. ��!ő�0Q�69Oz�M��.5!� ϨX��
����/���=�:�n�I�ɹ�-���3;ڣ)����8^��lX[�p�&�6P��^A�)�|V%�C��*��R.Jz}FSV����Z�E�%(*y`�)�w�@�v��gPݗ]axX&lq}�t�
��d�͉��N�ت��0�.�K�T��cB���D�G��S0V��1,H��;�B+���eCX�@���%q+��c�'�4��u>>D\�������s���5��۔;�t��-e��ߵ���~���l�>��S2#����e�]��k�l���NB���\��v��4��5���#f���ey�cO�=g�s�2���=Ay�T�Э�����mSցε}ZZ���mb����TC���I�o�7RJxI�4��+�
A��Q�����
��J�C�=�^�l���&�o�n�C��¥�����s��&��L9~K��z��3�ل�Ջ��:���x�,F�t���q�u��aUvsm����Gh�'z8�i�,��W=:Ppɞ:�ս�Ҋm5�Lg����������IwQQ��
~Ev��F�B�X��9T�������j�_)���D�#0�CV�U����T�P~*�jP/�9��{0���;�R�`$��o���㵯.���H[H�#����EĽ$Վ_^��d���4GԈ��4.�EI���7� ��Ri�u��Z�f��ԭ]-��"U���2�U0��d!#ԛ�Q$��!����7O�wٖ�gZՏ�j��K�����V�cj�*��F��z��n� `#~�S����E�>f�̕
�xݦ?�<�PW3�ɻ#����,�5܀�����A�%�L�X>���g6�H�k�C�H���k:�����74@�0i�O���O��(|}�O4&�I�>�z��-��\ KV�^���ǲ�u�v_4\�Y`޺!����0F��I�w���_��Y�E����t�-&��S(?�>Ӌ|�޷�at�'|��Z�	�̫�\��c���o�$c�?��𦩬�@ �l��{7�g0���Z�M��L�p0��*�,��L�I���$V�����S�bt؜���O��~���O��|�J (��!ކ�C=��Θ�3+/���.���e9k��N(���JG��㕇l��[M�_Ϩ��R���5rLe��Oaqj����P�A�+w�r�;�9�]fp�S��٨��?=���׎����)��;���oٵ��Y���j�F$����\ֶ���"��H����?b� v���P���G��A5��������,q��Hrd())
�"'���6�S{��<cD yUw�?��2��V?�Fp;9
��u�Vx�p��Ao�A���WS���iXl�r����%�V?%��r�Iv�Շr�̊B)g���S�x�gq�5tJ����Ec���=��SgM��m��� ��F���8f��e,��>rr���I����#K8��f��6!�a��ʛB��ʀI��,&���4x�Т�R��.�͹	�� BN(�3Y�������"�%MZ����pM��8���-��=�y&8b�d��N�\����X���?�ơг���W��.�޼`�n��WE4J~��/��mϱ�uy:� G��O���BHG�D>wQ��	iS�;hү����e�}/���jxh�X���٤���ҭz��oEl������6�&'�_`Ab�X��K��6�Ylc��Q�T�I�t���}NA#���?�Fқ�s�I�`�
x�S�H|�c���}���L_|X������n�3�F�/���FQi��D��xxH�4� $���A	a��V�2H_��������?�}	�� �X~�v��5�s�s �+�J�Cκ�@y��Za_FmQœ�� 7�zG'v��=t�\�(�����5�?�0�=�) H�v1u2�h�v� #�%@n�&%�c�����tX.߈�p���/-*F����2���|�4����i�<;����(�o��^�Q�H�}1m����8e'� ��ƼU ���_�Cj������vI;v�#Pcs��>_ZIΠ&�!���ʪ�A�P�O6�;�Օն}�+P%�l��M�#�X�ڙ�S�ؿ�*KQ�Z����dTARh6.��x%�ſ��X��������"24��7o�g�O�q�M�׿��G}��1u�<�Ns-v8�:c�{n��9,8���xn]�H))�5�ю���uB!>,���������TJ*p}� ��b��J�д�t���$j֜�1�5���rHEf�J�]|z�p�Ƹu���S�@CN�<�{_!�~}Z\�hу�NJ���.
��n�ߗ�4:-�U��ᚯ�g��x�I��5r�M�PK�b Mp&��K�B19��M'��ݑ٘V���:.4���g+6�LF'�c���R�������(R6�7���:W�q�>�>ܱ�*k/�Qq^�+e��?�����N���K;l�#W�jO���-|T|�L�Pd�M�s��x,>vt��M/.3���Z�i����V<�7��>�A�5���Fn�T3qj��rf5�Z��&���_�m�IK��^G�CaX��5�r�ٰ�n��Re��C���(�`���[��{�������sZ�(�q��jqEѧBM���p$@��(��ICa���G�[���9�Zp�x-�"��e~��<�p�ꞔd�S�8�S�U<xKCP�|;���;�����=S�u ���dBV"s�� �"?��/(��r�\�h�ǻ���n��#������R%���݃�U�Q������?�N?-��h$�h��s��ῷ#Q�5A'���5T�Oq06W�p�20>�)D��hn��p�}�w��'�S[s8q��&g����W����m�P�t�)IG6�p�|]��`Q%\�8���r%�3�o�jj)[�8b�5☸f��=�n!�&�x(
�Ժ����&}e�$_"�l�3�d.�Z����)p���ͺ�"�V���d�{�W��1(`�'N]���oV����G�Ka8}���h����`8�߉%��ғ�<K�'P��s�mf�i�.��W�����c����|A�-+�숕�t�D�<c���f����Ш�ă�����~ngI�!+Y׿I}IZE�.��B$97�1����z�I{8"�t���_�
�����X֮²*�.��i�2y7�ҧp(9!Ԕ\q+�7��e�[�'�鿳2��E�Sn��s�[���ݙ���oq�5����t���3V$W�#�4�u��,4��\�,ļi�N]�	����gU��� f�4�椒r�9��mߣ3L�l>�8]�5%YU|t�����r?��RW�����l���F\iu����r'������<h�h`|�ao���4Y�vD˟�V��>md�.fD��D����_��iE��⤹��]��˜��c�hL�g����c�&yy� ���P,�T4�X�RG�U,�TB�$h�vl2���P4�T֯���~m}�ىz_���'�w�0HZ�}���s����ͥ����ˊԷ��Խ�	H�mxd���I�D+��_��C�8V�F��#�(��M�.ᗆ��G	���?�֋}�`����a7eˡ�>&���\x�CG������Q����{;���6�#�@ؘ������i,	<74��Ut/��
t��3�6L�#��,�o>�Y��9��I�^ԧ	D��+�i��������7Z���||6�5!$G*+�����)�>4*�U��ﮒ7 .��Fo�yڂ����2��`8
�X��dy�he�ݟ��3�K{XvYI9�@��ү��4`�ҬM�i��gK
Y�\�
7���>�+6QLQq��]�c�${�O�8AL���F��i�:�RM�1��
�����O�$l��I�=)-"H����O�C����ϼ����|$+L ��ޒ�XPL��b'T	d&�	�L滫�S_<x wTG��Y�����/�V����W�jZ���#ߩ�}l�h�@��.��;�Y�]��Cu\�>������Z+֩ki�#�k�|�J:�<"V
B@��>*�[4������G���2����F��7�����68��x슥�	J�r�p��]�M�\{ϴ�o�FT]
�������*4���I��^1�,�[�I�����Q��֜�#�OՂ�uaF%Χ���ʛ�j~��i+�d�Ji��1�E�8}�<���r�����bJ#͋~��u��B��,n���?���Ƙ�e�us��������C��������oVn_Jv���&Ǯ�.6E�qB�a�qh쿝Br��pm �Ff��ݸ3��#u{{�˷�b!��.f�e��Gf0��G�Ϡ�*�r.���IX�A�!��X�T|�i_�vk�Af�Q�y���5��{��o���c���3Z���V3ڍ���m=k���7�ɣ�E�U�I\!K���'�hgΎm�T<1�$5V �x#@����T�7��	)C_��O��s������>�KP7jr�^�Ӏ�},����ł�W@�I6�T\7fZ�,����i9�D8'cu+�0 �)�� �۩T��\DTFM��!�z���'۱J�9�`��MؐT����w$qW��AHݠ�9\)Y�����D��]O�ȧ�ޤK�q��c7�Ĉ���`���sŰ�Lό���ݹ�����63���!�'�(��C��D���cn�H�}�T�J�h*"h�f%�w �C
���l����rM�V~����Y���O�gN���#�i���1�})Iy�C�TsE	}�z�������Ś��,�*,��d��i���w�����p�� ��1r���=�j7�!S���s���vÛ�Fh"Kы�v������L�5d��L(tC@J�9[t�"��-��{�������uP��~�	�2��P�g:���Lp^ֆ�(��0O�o���o#"��)�5�0��Y��x{f�ݔ�T��>�@W˙׳�`���I臵��C{�-¦����t����\�Ռ#X���9��r�z���y%����ж���-3&W[�n�a5�,��y���\��d-�L����u]r*V	���>	�}-��g#��`�QX� r��s.fY�ܴ��'%�o������� ��4���d�9\�	�F\d˼ ��O9n�ɥ�"���CZ��JxK6���i��L��-���)br24)��nJ��+PL;���-�\��i�Y�P\�O��n�16��p!�箌S������5����c���`����i}�ܩ�Pu�e���F_F.���X-gP�Bc҂A�K!�M��5{50�p����5N���}��^/(�Z��(���A���A*�_�9L�O[�[���&o$
3��d�*˫ky����`��~���u%c���n�'\&vw��,��\c���Q��V� 7^�^�����&�о{�{��@n�R�ω 71�O|{���+��!%s�K�V��P�h��ɳ�BaO �>��8N=�<��9��ϛEX�$��g�:u�L�1o�[�{JD�sL�Y N��_V`���e
i�HU�IO�څH�q�k��%�OU�}�J�|��[X��m�2���q��=h����Ĝ�<�ky[��hO��1Ö�|b�o�pCJ��?W��_
;�v#�Ȩ��_��$c���c�Lq��ˈ���7�?�NAx6�d�5�>����o�h�\�E��Z�C��W�{�*x��.�w��iΑ+�jy%��]�P��ƛ֫mzA�'�P�^grB����M�h�}���-&T�^&П�R���)�A"��n�|�cڗq�b����p�	r,���|8�TL<�c���0��e0X��O��<Z>:Q�(��ܸ�*Yq�t�wɪ��3x/s?(2),m�d�}dq�M���L.��'?���6���`�[Y!��/.A�3*u;\�_�iW�%��b�+�y���qy@��{�#�s*̠s�J�ά��G�I'��(:��Gd{���O��|���tѼCRa�7wXo�n��Xșa���5�Pha縓ʯ���>�4f��r��~���c��#"�i�i��}�o��n��3��T[����{K��<��	��#�¤��]P?����ߙ�V�[SQɖ����9(/�ċ[�x:c�Z�Q�{�Ig�z��h�f}
�GU����;9Ë$>$g�膟/��}���_k�,�RO����r\BO3;��Pr�^i^	1�?`EH���嫬�)��_9�?I�li�H�N]]e����|1 ���?׾,!(�@�-
[	7�} Psq� �J�Ѳ#JMTԕ�r�
PZ�F�(�T!��u���u�����(�C�k�:����s����������E-z�Z�&��zPHqRS,e�E%>���H���*���下x���M<��n�� �!�	s4"
�����3g�����,��r��:t�>��ºZ|��D�b`�*ݥs���
!DXs7�̥�����G�fK�Y����>�>��5�S�;Zy�)S�2U�qS����ʬ�Nc�G��ӏ���_K�7����intR�2�!�&�x��6O������?��O���swP�<ve�1խ~�Ѝ�$�j�=ߥ45z�;��rPYSz_�%<yU~
��=�G��]��� �"���i{EpCR�,�q��Kk���!�@����� �����jK�"k Ďv|`1	���Ik��U6�h��K���sړGu`:D��qh� ���UQ2A�����^�lHu\���迗Aӧ}*b��˕���-�?�	&��t���=�	5�� �$<tj@]t��Zk\%����*�1jM� ��_���o�3�1v���B�	�7�r��v@�Yv�j��r���q�0����Tm��cQ$D��L�GW�>#��K#�6_y J����G>�F���ߏ0f0_h͈���,k�����Ŕ�FFrHPf��g��;1�c��]g�����Ł����v5�����)�)�Ҟ��5���ԡ�����	���5`T
]��v����5�=}ߥAyʖ��E�J��ik�;!��-�q���ue�I��r�L����A�j�Ŧ�8�/'��$�G�~�e�(-���k�֑!�[/j�韚�����L;
ycq��`��4ux�?�<��u��?q�oKB��n|�E���~ɍp���1o 2Iqm�:X��Y,!�&a�Յ:k߮sH��8d������1���U��s�PN��X4��L�-��+g?��м)�E}����7zE��g�``Sw�6$w9������iҢ6�t~���"��Ǹ�#�f������>r��wZ�_���%a{�[��k�m}��'��r�#$4:�	�D���B8�*~��.�s������I1>&J����="�Tj�A
�k�#��-7�G�\�O����!����k�#4��3�-��Ŝ �
�m?��,���ߕ�Y��`t׍M���CS������T�Nn��\EjH	.".i��nd��Ż@/�ľ��SG���)�G�_F��%�؏.Z���*�ԉ_�*d\���1����(���'�?���B�J�SK��\;^�"*1Y4�WS������?�c�� C�j��a���]�̾
�v��W�Qc.�B�9vuq=�{k6�>b69z$ϯ��Ê��&����S��b�$��x���7��{���ﰋ���
�ֿ;dU�Els��HtvΚ�}t��SB�(X=�E�ڜݞ�g_���k���-$��T�/AV��'u���3�W@��m�m����]�s*����L~}*6�Q�^����Ϭ�e零D*�!8*��u�]nAig�!�d]9��wZ�0ΙbrHL�M��m��w�ڠ3���*G�@G�)n��ۊ����u�t�K�u�7��,�Kf(���Q|P7��$��h�2b��ס��V]����әM�Hv�b5�U9� ^F�T��Z��j��JscV�kC�_�y_��6_�Wlx.qT�?���3��=打�g1�m
c�BD웲�^�~r��dNꡑ"Qu�A���lo��1����&��T]^}W�v-=�X��c���t�T͇�J�A��rZ���Q�Ϲ���h��R�;-�cfW ދ\�|g$RZF��X�g���Mh�vP"yh�v���}k��B�'+�P�H��zP��',0��^�vt���SkTZa�/=S<��a�L��� ͊�w����)��?Х(B�L�h�X�1�T�) iO�V�7Y�C�"����0Bѩ'1��|�*�o�&wZ�Y�'+�Ȃc=Sk���_�
����-���>�EU��N�C9�V���3�L���Q|��!p�S�0;f2Ŕ�.IL�����]{Zd��g��wD���`zn�9�*<*��n@8����UP�[iJ��G؁�v
�JԠ"��f�.��-� ��h;������N��g�O�t�sk�R�|��^h�&���Nļ�Sj��^�+jZa��%%��W�H�ɾ
�|7�=������C�:���QL��D	�e^��<�V8Lgh�������`�Q��JL�S�@����w�1�q��;<�9��!L��JK���b��j];��w1�t;��
*H�)�"6�-G�8����õ7��-�}(%�^����&����W�����7���ӓ��l�M�#yЂ��?�y�(�+�5,֞<�PΑ��2�n���;W�	�TMH~d,M�|ղ{E��į�W_����z5����\��g��U��l��?�_�h�@P���uL��(ַ3Q�U��%8����2VP�eu��ڐpj����A~,��������pǋ��h�"�0�*"�бFp��:e`=H���E�VQ�'���$�ɓǜ$�za����H����(�erVy��n{��Eh�U�������i����ᅸ�K�R6J�+q�^#m������B�5g�w�۶N�G^u_^:�h0�C��Qs�D�q�v�τ�͂qp���T��d�o�La�B �=�F�3Os��q���f��\*�1	Biɽ���!?>u��ɨ-��r�O]�4�e���%G+����^�IUG�U϶/�BԵM��.s�mIz���:�/b�%���)�z����rBt��0�x�a%���n@F�N=�*�Ծv�(��H�y��P]~��_X�#
[~�b����*�l�uH�W%ɠ��Y3�S
�#=���giw�\�c�m���������i>q�n���劏��F���8��|�"�r�����䮕F$L�u7��O���d��k�0�vn��Byi�5��J�4V���7լqc���ݹ�_2�=D���:͔���΁��T����ǻ,�ޤn0i��H������'�BېH3�ݪ��߿:	P��Rﴐ@��'IB����jmp��k���4�S�=0��{?|%�
S�sZ��3��v�Ϊ�o�Υ�W|�z�9+�]�R��,
�]	3Ǘ��<
�%����̡#���r2��LG����6b"���еb�}\y�x�'@s=_`�~_�X��%������ycΥ=��$��a�BOmom�0�	j6�8ev�^$�4J+W�e8�@�M�)�
��~=����O�a�3ᴞ�kW����={]����QV��"ě�,iC�=���m,=H�${��f2; ^hD�q3���r�3ő��rxz�0{AM����g)O�	F�is�h U�H��ع�u+��X�����'��@͘^�X���g�,�.8�<C;>���*`��a1��];����y,S�/���{Ch4�,���Ǉ��h+i!n\'�޽��e-h�;z��}���3�bmv��.���fc��웆$�o��Myw�d5f{�F��<,�9�y��d�K�g�)u�m��i��^�0�lkE�e��y_��)�K��/\1�CR��av(���!���Ng���r����M�P�w�]�V�xo}�0�]�ZՍUnk�k6�G�/B�*z�jq-�l�/C�F>��Q�D�}�I�u"V������5p�̖^"39Ȭ�N��N�NB�nQ{N��n��H>�����dg� *͡^�I1�J�ƩT;��?X�٥*�<�S�Ww!5D�V�� 'T��D�
�