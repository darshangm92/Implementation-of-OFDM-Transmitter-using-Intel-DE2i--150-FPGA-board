��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<������M�&ӗ. ( ��:���n�$��j/N4����Y���;�{��p���&z��>-���Ν�A���E��&�;P��1qqzf����H<�����C� Vޕ���߆)��ڊ�U���|� ��_:5	���cx���,c%V�թ���k=�U4���8ߦƤ�k(���5
���5�$A1`	�NU�˂8[,D\�3=I���偁WG�	/��`�3��<��W�2moڡX��S�1�d�Cg�~H��E�b�U�d�Lϴa��]� ̈́�ڥ��9#i��К|}3��CSk��P��O3����}H$+�q �p�͊q�k�K..rQq_>yE���0�����X��W�Cӕ��R����̳�@5��m��_ZXJC=l���wTP��I������d$Ã�c��D�_s�'��<F��}>\dK��;����������HUU��,* j��ZU��5<w����lm��5�t���!s
1�!�Yɧok�:�$�>�w�|��1TLVCG��b��1u��c���ANT�疰� P}xOs��+����0t�R]��+y����]8��D�Ċ��=4��4^7�� h�����Yir�B&��AJ;m�Ov�Y�M���!�U�8x�'��K�М�7�m�X�JVi��X��n����H��WC3?���nk$���:��[���H�gH�RRK_p�듭������eD�I}z��bm8[0~�+<�;�s>E�-cD��u"�nҴ	�!�n�W1� 8+ I���Xd�D���9��sW<�a���uӐ�HK��*l��A�t&n��4/��7�e��V'�9�*�[t` {�|E5Ј�d�q���a-p
�d��Bq��3OHo�3�e�� {������5�@�1�Pt�K�	CiZ���{n���Z��d=��u�>q�0W���*�-J���i�t(K<�9s����H<�h�ה��ȑCC��Q�lE^��N�Fl�kLd�O78�3�׭�͖م����5����i����g��:�\�b�f~��aMλ��ϯ��UN$�9�cI)��v�ˏ��d�p�����w����F���E�=f�N.K�X���|ѹ�^� &�6�����Z�}�bf�́e�X�R��w�>�|����q��c	=������	�����~$Ō=I�uf�!�V���T�N��\��	߰�9��?�8��Y�<;$�8T7�<��G��!<��6��~]2�~�2 ��p��\p��]a�m�-C��M�\�c���χ`�k�8�m��ݷ��Ӄe$�Y�#�+�[�2Ȁײ,�-�n��I!ױ� �&s�;1���u��EĀ��E��4}@͏>U�P�C�L��𴮑V79<WM� ��f��4�n���D�*q_e��Is�1��*�g	s�O��4
�c��:*�ٕ?��o߈ԩ��7�ݙ����`Ű3�){�hR�)�`w,؈(�R>E��)�[z&ք)=�ɏ��ql"&��X�[���-Mip?���%�}��㑝�H�U	����G�\�S�M|p��F�U@d�8Ț�N`���/�l>v!�D��R6k�X�y�^�s�6zbr������+����F���95����Y�$����dq�eZO�	��f6�;nm-+�<;���u\���6?�)���W��Di1�U�E/�+]'������q'��˫$���9�]Q�[�xپ{赤�AVb!U���؀�[�Vܐ�7�T�n�{#��.��)�
۪�`�H6��w���?�*��70��� F�m�~�2�꾒B��i��
!�r��n;�(�ܓ�Av!U R�-C���TjJz���6��%����=�O*k�
�����4�ԑ-�N�)�S�va+�r@>�4��&'��`	�����-B9�(䳨ܖإ�G���ѡ�	goɸ�B�Ed��\n�>H�_���bJ$�G�#��mH��JX!�u�4qau��4���R��Σ���]�z5�W8��҆$	� lSF=m�h���Q\�
x,�[C��"�y��� v���0��Id5֒7Y��X��H��������P½�ZK1�wP�j2�>����P��r���F�S�H`j�͉�w�kO���8!t2?�+n��YX�{>ax=���T�n_��手$ť����j�to��s�(�#X�Q������Ca�ASϤ��OU���n���E�t��0a��⽪5hY=u�TcMQ��=�~r���}��e�#�,X���\�ؾd�D޵io���xP��.�b�	�L������b�|3,T���i'	��t�2ep����hS����\;�ZG*~j���=Wg�+�{���yM�JX2D4sMF�Xcx���h��)}M��<��o�J��g�*��-�����{��Ll�� ����1.P�=�	 �~�i�.�-�-dC��vr �4�5��yX$1�t�*F�֛4��j$́�ʥZ�x���#T�f�W�B�\�"J���JEi�QU���6[��y�N��Q;�r�ib���8�F��o�s�\���9������t
��b���}��|x�7؀)6��p�f�JꚄ)0.�L}�9��O�����hjNTS\��=��21��	gl�詀���:BOr<;��͛>ӶB<5��71�����>j�oY�3If 0��KF�.�y;�Z&������c̨t�)4�F��a ���7���h�KI?��ߊ>�����t���N�\�n�w<	���
�V�#��t�js,?/���,��~���ru�=6�ޘ#����(��8�U�lG܅.��K�J�o1�X� �n2.���8V�9m��w
4�yVJ;�0g,�G/�$�g ml�Ǘb��×)����H��	�U%�y�����i���\Ю ���0��]1��xt���[U�
](A�֦E�zfd�ulY��f�]��\$c^c��0���[�Z�ˠⴙi_��+{�m�A���mH�8"���pW.���[<e�͂��M_�:��S�t^�{QKq�K�����;�pfky�y��B�g�^|\i۠�������Β5�� �:5r�ۯ_���2?8w�)�t�ʤ#B��������Q]h�4����n��瀪�4�R��5	�Y���(X��S�/�s�k<�yw��85Yf� �mG�f��f#�=%�f��pU���p�Z2c���pk�xҠFh����x0�6��:[3��T��!�9���|��1�i�H1����lpt9���oI0����1}�2&F����M���#��e�w�)�I��K�V�/�s�p⑖s�����zʣ��]`��tK>l'� <���x,4��5E���E%>�LyI�0u�C����P���r�
d�.�
х�!�lWG+I�{�<s>OE4��3v��VՕ<�?�A�`�aq���`ۋK
�>sr�.�x����9�_k��t뾗�L��=��zVn��S~���	�{��Ac�
8;���|Yt� �����סst�O� ,we�� OX��b�<��B�=������B�3��x���^S��4��K���(>�z4jvlOO�E���2������l���%���j�z^A�q��#3h�	P�J� #ll��q��0g���Gn�s�I���ݺӶDE�R6ܩ�ػ������RS,֑6C[�'e^
/�oL��"*�w���³ ��qB�b���T~�;����l���`��5%�`$:H凤JJ$�|Y[jt�7s�B/0{ ���]Lh!Q,1
8��BƫN�=*:ί>٠!��}Fx�b�P/����Vg�b[aSE8s<����D\�;�To?�@�=t�*�+��c�ή�<��u��hc�;]9����v�`���"Jo=���؅��c]�/�͇܃V�����}k�eΓ���g.Z�oW�z��[�v�e�)@P��VC���s�J~�,��.^�j��2�>�ZK��̎�I��8���Ѥ��0�ԃ�l:���#ø3qWCR������A���c�S��G����|�
�H2֨�5�gJ�"�b�񧧑�(54(�T� �%Rx��+D�'�08�f�Eu��~ڄ�<�//�tB���L"�	�f4���I	��ت�����i'M�'D�b��'������T���a��F<��A�!�e��j�sϬ������Dv�uY��t�4�� ϗh�� �I3T6�TJ@��� P�,_�Ɗ�u�����7��ǚC��Wk�EK�͂;6*O�{�@�F ��Ք�J�4��;���>�R��?�Z]݁�y�L��$K�'L٫��ڦ���-Mu��	yY@�z��N���ҫJ,�cɍ����ɵEb����,6����ns�����7`�6A�Y�����F�lU���ˋn�u�R�&c;���
�I�=/N[�n�I����@%`�R��%j>4�R僩�wP+�Q�F|���Y0�4<t�i�j(s6�'[A��Ĺ���}���r�o���v[��&�kQ��V����].%��� ���\�����;s�.�V*i����Y|�Ndhm90�1 �t��V��OT�p�4�$x,Y�?�e�PX|5s� �Ț�ϸ�S� �q��v�8��3-nIZ.k���=<G���RӈX����ߛ�SE��iWb���s�ZiuD	yc����4T!�.S%_�����������H�@�/#�3M~�#	�$�ں=��������L��4]+��B�(y��࣢0��r ��̦�L��P��Ah�(����G��Q��zj�_�T7����v�5\�d��ƥ���O;�Ё\F�kB|�l1��θ!LhO��4Q9��3�(H�{�X/b���C�<��WA��i��wd��<�ѻ3kx(sH
Lc� `�&�����=9����6I��6�c©HOԝ`��yrYƬ
�5��|�z�w�QK��W�s���C��[u�����1�˝�lCP��O)Dz��k�+�Yލ��r������!�����֋�!�K��Z� ��(�tSw-���"):���&�~�.2|&�f�$B9Ū�����p�\��e��m,� k����Е�7��J�]h&C=�š��C�k�.���=�L��!o)��Jv�vE{zK=5��/k����ڸ'/��̋O�K���z���7 ��2��gt��sӶ�S������N9��&�آ�|�^5"�ԙ�|c_r������MFA, §�P!$�C3���Z�Oub���K�5$A