��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�/Fw��x��b ayk��]���
t����jw-V��k�d<a�f��xx�/�~���)ҁ�چP�^4�#�Hy��9�=���
}na����ʟg��������lE�R�6By��������"'Zw����k��=y��9XmLjp�՘`/��z5 ��r8���˂}���\c���ô5�������d<�,�
�����f��t�Ȕw1���a��Eg�z�*��Ùk��W�[\�]�Gٿ4�@&Q[�t�&8�$���-�PC�����M]�����9���4tT���Y�\~��Qd6�ݼ�[0m<=R�  �@���d��}.lP��+��=,��:�1�M�hU�c�[�������<��m�?��O��Q\r�&���c�Z"f����1ox�v���yA��724c�7Bb6H�k��e/ʛ����(kvq�ˡVK%`��We &g������)|�|�������o�7� =�b ��8��bLc~�6|����ݘ��JC�E��m���+پ%-('�@��|�Ԉ	���-�P�~铛3$ӂ��j�ص����(Wp50�vǽ�8�o����gKOz�鎔�&nS&X�<{�Ҿb�>��s@���}.�:��t,ּ��~�cMl�{�)^�����P���,6�_����6����-Y� �S36�nO��DZ����ҋ��`�?�͇-��T�
�fS�Q!-ض8���=����-@�9�l����~Ȳ�\}�=-L�KQa�f�܋LK���}��\K��n�`�ԯ��WT�!��$k���]_!�׫t9f�� ;Pq��?�B���; �X��7z������f ��.��� �x)��m/%>Ә.G�c	 Tq@�v@{��n1R����q~CI�)�Ā�/߂@��w:2���dވ�V��%@��P�}DV�1����݈�:hs���l��J�����L)���`��WmS_[�v�L�O^e��X��=�����,h��Կ�o���r�����D����� I�v(�j|2��d}���8쒝���_�r<he(��L _����Y+N@��dО���4~������0eMf�!B��MQ �P]�Ó]����{J��M����C���_�A~)�����i�C��x��O�������w��9�鳎�ρu�\bj��t<�B�G������B�g�(��K2D�q���1Q��(c�)j21�E'�_;�	E
��Ik�������n̍Iї��"c��Թ	��G	��yq"}:E�A!���?���4��m��hh7l۳�2�yܓ�M=�j��e�(Q���p�	�{E�9�q����霰�$�����гp�j��B'9�@�n������{|�G�.08�@MUeiu�e���,��1+me�Itٰ&�5��P7�� �@Ϝ�c
�?�2w����
Y��p��w��9Z+�s�]bң�iH��h�`��<�͂����wU|s�=�\�R�CJ`���(bKy]�\�%���Z���.���0�J���1��]����OR�v�֥ a|$�{��iW 99fZ�h���o����H�w��xj��֚���$��7D	,JAm�*�/�}Kڶ�ʁ��iJ�p�'�f^Q)����x��-*e	B��l�����m����`qf�Z�����P�υ,7�<��rD�԰���\W�Tע�����Gz�Pԡ�'W%15�{[ɷZ�R"d3���$�'��S����Dh돣}�����ln������)9�D�9�y) ����]|��9(���3!�n�]�c�:��g�����}l��L�%a�d,gf�W�(^��Ъ>�'�Ϸ%��ƴ6F��F�A��)�9�B��uM��#���@��C/筡F��.�πCy�Ys=���r�T�J:�,��3c^RS���%�l��q�#a���|���:��,��I�c��-UB�P���y������g�g�!w`�v{��f���80��6>�x�=�*�X:N�!��i4ޏ, >����r�Z5(��p�v�y��EC��n�[g`����Y��e�X��u��DM8��$N�D���6A8}+��c7�)Z�]�&�%���j�@{VlF�[V:#��)遲D����U%��|΄� ���/�����-.n�p�3UY�,��@??�b��s;_n;ʫ�:y�
.��0�N�۬�