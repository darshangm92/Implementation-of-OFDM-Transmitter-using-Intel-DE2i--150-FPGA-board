��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����{�sGq�*MO,.���buD�"���`aő<��<XB�:K�z�9�e~l�9L0n�;��a��$F���8{�u_٬DWdZ�X��2`C��o>r�,��<oU�3Mx���C.X�,o���#2�`Z���}#�9[�{������d:��`S�޶e�s����=��T8�X����܌%��ˆ͒�E6^�Z祈3�n%b��_����x���A_oWt���)����.���[q�p�B��;�����ey�s?��#�ﲪ���ߵ��ƭ�gl��Z툪.jϒu�i�-�*�(ދ�AT�dM=��
\��l��i��~�[I�<^���be���^���y%�&mL-�*��R�eAħO
��-\���$����\ڊ�v�M� �!���E�\�V 9"J䀉�sl���$w��4����"�ߗ`݊T�ȕ���"g����J$ʀ��v�ux���4�xL�K���G�S��,��XI����$�xd=a�eM��x_�;K��t��)� ��B������HT���.Ů�)w/�:��9�����a���<B�.�ǸѬ����/�����/�-y�Y�&������޻�Am�\-���;�'���4y�"�4�4�N�7rSKv%y�g{tv��緰ɞ��[�ȹ���Ů�ñl�YӤ��ᰋ�na�NASU�`�g(���32�^!�o��c��0���=uk�L��ƽV�b�CXI��:Mz�����I��}�����*��`�~��İ�  B慜��HJ���
�i�nB��Z$�[$g���7���S�
x~2Α��Ƥ�F_j�7�����t� �	xD�,ȵF��IG5/�&���Jt�����2� �����[��%�|�NՎ`֤��A��/�����@��9���#T��fh�`�p6v2LE+rY (�1<bS{�T��(����a�56N�Ӫ/4�SE�fS-�=�Aӱ@@�+o��o��N9)6�RY{JB���
K�����בA�1a�=�hM����;!�(��(�<�57t¹�o�)HK�!�|	YTU|�?-T�W=%�;�7D��]���1�4�cn�A�q�&����������Bg��]D���g�~��m���!A������ˀWYɞ��<� ��T6G%UHe+������'�SŘ���쳆�x�q4�rD$�m7�1�?�]҉�o����l���5!���g�/}�I�&w@[} ��['ҙ
�/`�ka�;c��8���l�yb��y��"�eI5�G��K�R��T���D�JЇ��"�Ĭ�p����U�S�;�4���'�s˞*τ���|OnD�="[�	�<�]j�iⵣ��j\|"�$�&���]x��Z���j|J�i22�ѽ��y�O%��\\���0o&"$�C�)������[�=���A��s,��j<�Y���$5#'w��^b�
6��(fs
ͻ`.���D������M�-�9U���%C�/�÷�R�I�����81I��3���e��ơ_�V�Sߺj�6��}}� ����%��ߓ�znE�Q�S嬛n�����h+J2ų�y��C��~����(cc+Hz˔B�]�G��癪�Wt��0+n	H��=[��u3�9@�'�jvYP��GI�o�������fr���F���<�t���d��+��	<Ș���א��,$��ky�^��0S��]����
�7З	��w�O
]�8-څ��o��Wy� |��?g��Gh��������xT��ʣi�2{'�WK�UI�W3�wd�]�&e>�t�'t�Q�E��yɅ��"��2�dɓ�_SP唈I��~C�q�i=���o�c7�;paR5.@f#��0Kl��V8ڪpq�کɉ�R9���U��޴p������LQ6@{�G>=?1�T>��:���YTc�'�U ��_-�<�p� R�^��I*?�ۡ�i����H�Ŷ�%���O=\�Ȑ�k�,��v�������㳀�Ύ4J�^�|������B����Z��}�ͯ��/xT,U٠�r(:ƴ���{Х�@��8�}*��8���Ւ�,Q�t�y�6�|8Ѫv�-�����힨����UI�X�.��U�il6��F=W����M�̙i"�/���vv+ު�|�p!3�| ���i9zy�6�����Y�ˑv��X��M�, Pµ+:	-j��q��I�ӥJF��nyV�N?*��8�J��)΍D�\�+ZJB�Ŧ�����>�þ�r�?�!d՗u����[|j�=������L�xaK�v�M4��۪�L_��xpa;�z��u�W�LՃ]�=13���{��@iى���%�B�I�R�#n�������F���㸉�%�/�"-�	}%Tާx��:Ը�0�wd���Y�o�m�)��&+W�T����� �=��piGSԴQi��;}��s��ȿ1����5�ݑР��e�H�Q�Dʛ��-���^J�9$��n��w�_m�(wq�ƓWih��7m�P˩�4���"� 굄���XV�����6������:�X�����(A�/��R|8![�m�ύ[�a�.�
��&�z-�m����(�5һ4e��<u��$�۬Ҕ?��=�[�8�t�P�i�?�t��*U�J3�j���o�潦z�OL;��	H6ZO�i������f��i�;lZ�&m���B�{J�q,Y����-�k{ԣT� IMإfPSy�L HӠ��'����?s��t�c���xE�^G���+�̦�,o[��ȇӈ^�*>X�p�H1��O�c���1��㧧�%RS�,w�y��w-��N�=����-K
����`J�kob�ϧ0I�R�'��tx3.���ޕ�&&|t����{18�|���L�����R9���A W��J��<���K��\�hK�֣�ڕ��4;m�� ^�&\��S�S;�pcEE�%��h= d'`1�99Z�ތ!�|C-���)jt��nVq�����-C�R� �lXG`�?�qB5���J�F�.ԸK��ˈ�g��@�3����!R�i�>��Z�7K�Օ����iK+�Χ�ɗ�������*�Z?�!�|����W�j�i.��t}(�S�����a�ȴ"���P,���l��@M��?�>E�y��qKDi7���(��Y_T\��CTx�c�~Z���#u3aR�h��z���)�ԗ��q��6sM���?�6󻦶䱿VϚ_
�9�Q�lPA�w�#�2��X�Z�f	��K�׊W]�WԙmKc	�S Yq��Q����ɣ�Kf��*����o}�y+S�[���
93�얶���lW�-�zR��� D�)?}�2��I��;�
U�l@��uck���;����t^�m�����d��IO����n.Aw�F{�y)���i1����}\�`�ø��2gƷ|k��k::!#'����������M���M"�`��k��y����H5vUQ�ѱ�!і�����
1��k��(�B���h��wW�����?��Ǫ~�0������f���N�H��h�}gPˋQxi��>�A�$�'l��{.��?�܅��_T�����i�7����༻�wRS��_���P_��~�_�AgZ|e�㷐(��t(�}ͩ�|#Ay�DtNJT�>aU�	K^"'Yj�dk2U���=B�O�K���aUOP�ȵ��J��:��gĎo���à��#4oAG���`x8��Dx���%�+]
�V	��a��55�