��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�RWG�a'hj�hD��h�\�\Ʌ=��R�^�} ��@��z9�|b�[m�X�7T_��s��'�m��#Ԧ�P�_B���������
�A�l�9{U�-�u�5+#������	b�J�A�`�6~ʁ*%�E(�x�:5��]z��j?*���GB�okI����"��zM$�&L�W������Pd��5����׆G�js��{Hl0(nR��U$�,��\H���yMO7�d������d9�52��f!H�"�k�R����u������T�_o���k�:$�'y�	J1 �i<H+����G�zWv�Q�PI�a��jXὠ���_z���u�&'��#��̛�3�
�)#p(2|T������"Æ�$��6��tn��0���7�%�D`�@���=�e�\���w�+���w�\[Ϳk��y���m$�@�ո/1W���;J��� �;I�h�?���8B9�X�,TTtg��3wR7v(�E���]z�H�B���1�ݶx��w�ٚA�6D���<H`�G�,�uM�mq����&e`��Ӊ�ĺ�x=���~����ӷ��7�g�|�\�9jD-T�@,��Ũy9�	���;�S����=�X�(�q
u�G��;䢛K)��&B�WE&���������C����O`�����8*�e���g���_�J{p�J�Q�<�3�{�T�d��W�8�)>� ��3�_������?K�����H�=jD]n��4� IE��΢&��I��D5;��bZ��a�1"{�s�l�Nd�/$��m�4yD��5�O�}4�:�	 ������9��1��@�F�@�^m=���1�g�+��l�ai2J%�wY�|�R��BNR)�N��� ����C�
zw��I�	gE��:�
���U�-q(���^��wK��Z��v59�T`_9���?�<��v��k au� M�n��|���8U�l]*�҃�*�{��퐵�̰%&�W�Y�R����#�  �k����*�n)�
����ٹ�Ӭ��2�Kgo�Q���OĴ���H�x���]n��m�(0{�PUwQ�b|B�L�L����֋Y�WJ�.�kɛ�)���rzK�|��q^?"O�$���t'O0[�2P���"2Y���Lk��jf�˼�kz�g���'T|�VgZmo�Y�a�8D�C,�7�E\�R�ƻ^'�`mL������+-��bz�+��f��ד��@�g����<kY"��lNH������p�\�������@e||:h(�`�	')Y呈^�Z� �����a��lj�H�6g$�c�E���`"	Kl�#:(s� [�(���3 &��_>�9O��z�?���!���7�|��M��SO�+la�r�R&#��s6s3[Lx�-m��Kep�7Ӷ�L�fx.2��-��	��7�E��zH�C�� |w
��V'��9�D~=F^`]�t��3�E'��̬g�F��P+0�%?�e��� �k�)�З�W�Z��r
٧�����fx�Pg�P�7n�d�'�Qԑ�zjR��$��:XBC���B�S$�Y���1�l�;�E���NO8cfS<bD�7ɯW<���C��:RF0���-<)^$
a�$f���S��Ca �����B�%��_����'��"�B9��=ň
���T���f��Q:����.�S�<+�	��
��d:�����Q&��������'��P�EcZ�)���N�$Sι�D'6j�eP7�\�
���/f:)�����]H7�Z�
�����]�l%�т�#�WL�3��'�]oq����$���T�@ʥ>�g�i���z���&u��I`���B�
�r,���He�	/`'!,��=�<�X���-:ˍ� M�"�ʥ=���5���&y��@ ��K��u����-�.��%O�~�J5�L|���5���ӛ�5m�P��~�0�1�3:{��z@�@�t��A��I/NMgqP�O���":%AN�h���Fɶl�<5�O1������/"�íˉ#3�ixKݨT��wV�0���Y*����������Q��`�Y�)G�+>�9�:4Z=8�n� y�e��tOI"��D��TQ{�E����(g��~
�e��F��"C���i�U�/h'�۴�l <���v^"w0��!8jG %��]n8���6u&�D�LlERU�J~c^e�c4���1�Iv[\C�ĚMM����@S�������%'�w��;���J��p��X�-s�D�Kx���l�]m��t�+"ȶ�7����� R��E�ֹjm�|���eo��'Ϙ��>��Zt-+��E(gy�% ^��3�8ƫ�~�{�A��o��KV���q�!^��6�,�r�|r��n~���K�����Դ 5�|8�Y:�E����*��|��
Ai��G���������������B�53��e�I���G�P�WLó<Q<�E�Hc'St;@�~����5ܗ����Cs��j�@�AY��8�^��Q�U�¢EQ��o��gW{Tv���+6n'PVHZ�Q��tJ�,�-�6m/M�h���:§�5�A��B�*\���0�|��#Kr! ��:����lF�J�*�YFy'�>ܢ���h��Nq�U>=G�>e������,�@Hw�,�S;���,�����j����u
mN�M�$���x@��<�;4���
�������.<���wH�<�y�����vӼ�gΜԤi6^�b��u��v���@E��0���~�"��%a�4vj�^��z�N{���#���ǆU�P=	$��$�eK*�#><=�L5 ��9�*9 f�(ˉD���l3X��
�|�͘�Z���s/�n6�,��7�����-c6���-��_�S�k��<��0'�0�����Q����~��A�TIe?s���,�!K�A�C	�X��6e94q�5�P9�Y���L�P'�H|�ӅX��N%'�&B�|�_ki��攦�-�>N=�;�7� ���c�tI�I����h��������@$�²�2k�Dl�H�g��jF���< v�j3k�lϽp��ҿ�2B�(��2��;�@`	MG�K�N������r������ń�P�訹4*)q��b�w@(q^�A�[A<kzZݖ���@�v�D!R�.R$�Q�K���d��1+���6�[�d�6��O�7����s<;j�
�M�Hة�MR���,+uv �;^w�NO����������?;?��Q�W7j���/�yG����a�4Ժ���~�����bA�V��f��8���e8�=w��̀n��;���5����m�n�t�(�i�����(�#1WH��5u�T�8(z"ȵm*s���v��MvL������ÓHv��z��N������Ь�؝�IpR�>i�Y�1-�����Iȇ�eW1���)�v����;��"=�6;+���4�C2�uV=�sd��Nvcȱ�{U�F���A��,���c��4���k�Fhh\�Z���}�d�U�q9{N��m�	Hk�u�o�t����`�͈l��\��u����4X�B��I@�H�ao�K�56�j�aS�`�<�Θ��x��#�tj:��������	��Y,�#�k|oc����Ұ�Lw�Û_U���� 4�u�z�;�#?�G�v�T��E�b�g�ڸl��	��[L<5������QH�6n�Zkɕ�E*P�,r��ƦB,��~�\}�u3�&MO���g��ϙظ��z�46��*T�?�y��دX�4RUamS"oW7(gE�c��8V{xG<���ky��G��ee�J�5ԍ�J_����1����\����}�*4��/�[��$�
�Ƈ���ԏ�<4a\��@М�ٷ���SS���Y-��}���',�}��I�>�@q�?OQ�Hm|�w ��^��� ��Y�L9'b��Y��>֖=�3�J����S`�{Vf�D)���D��+���-���m��.�����č.��3����&/q�7��5Y!.�<��8�][ �.�B��j�E������`���k�#`2[�]���5]���|��t{��x�x� H��]d�"��V�h!|CJ�3���%���=Dcu�7�8fuW]��� 橳�2𓣮vYd�WB�����;^v�c�4EiB��K�ŧx��ǽn�Z-��Q��g�`6w`hN+R'�3�	��4��h�ƞ����w���e�D�e��2RE`��^<��`�aX}ᮏ�z������ww~f4�
�\PHC�I�)�9���ސ[��q	Ɩ��w��*�3�2~&��,�wU��vO^�^S���:;덦�٣�t���$2�Llo�6�����gQo��֊���<���1~s\�T������Tƻa�ed���5��҉=�f�v�pW���ߤ'zqRȦUC���9'�>pe�Ȱ�vS73�15�x�����V�?�����i4 �[p���#(�M�*�onG�8�1M¸��9��ImOt��Ӏ�"!��F���lR��s (�Y&IǸ�BF��<��<�ɕ�<�W���n��DLJ�!��S�,Qk�pw��\ <�R<��9<���m�2x���`���:fr�i������Q&�N�N̉���(EU+�W��`o���:E\���U=� ��ΧP�pCf���`�'ܬG'���o���Ш'_A�Uv�����v};&l��'"4�wZAƐ��?Q6K�~���%�I�F�uӰC̸7esT3���$㱘��и�����F�;2��)�_�p�6q��i�:O͹r�<۩�z��������#��i��.���q�M4�5-s����Ay��*�og7��"����X-x�,���!�Mr~L��6wf�6�(��Ît�2JR��pי��0�����3m�y��]����^8��N荑�X�L��	W�̧	�l����Gm'"�i�1��$�0b�u��D��7x%����L5�����qH>%���mϮZ�@Gü�������]E�PA�>�� ��|��W�5�n��}�w��F�i�F�����WK�ԧ�|m5�b������o����#Y��1d����l���0��@�`�W�'���:�_� ��Ƅ��'4���l<j��j���<<�x^��S
juH�l�����G�I|�
�?�����{��sYߐ�K´�#�޳�'�x��]%o��ezy����z���ozA��B�0���T�wL��3�Cw�i�2����	 �� �tdcG�	R����`�~|�ÿ���fJ3�v��	1��L-J((�<S�]`�}�@���4-��kkh�f�IC���(@��:,��W4ev��+���iE�\�r�sSzf 
W�� NQ���gq��٫���E���[��vzT��3{ř��Vp��n��)>��D���z�� )��5�}؛��	��Źz����F>�Rλ�j�NZ�F'+ZR��N����j�t�e��Ir>Â��e1.�������9�֎/r���k0#��S�1�����H�ox��R����!�� zY�[ɗ�i6Q��li�Ns��?���O�\�Ȱ�.�.I�>�QхLz�H�`��K=�s?Z~C?��6Ұ����s_.q#�c�n�Y�]�z�9�/$$��-�\Y;�+Ā�tDg���/�P���Uӿ���*�$$�ٍL0a��.I����X��7M�7J*[z�˔+��3�j7����=Ƙ�ԉ��r���	�Z���|.:#��'h���vyi�%�HI���~���7�8��H�I�R��֨��i�\N��}<we����S�y��I��oX��VH���җl��Q[�X�]��Z'�Ge����b7f/
2K2��*U:$�9'��A/*1Yq5�����/fO��08����B0�s�>ބ����&x_κ2��T��َ����m_%���\��CS��d>��IM��-�[r�,+c�X@OD˘��H��6�]g@ş�ԣ����ǒTi�E����/l�i��b�z�8^q�@�hC��9a��uFÓz��0�Ǝ�܉��ۿO�a��&�;��7MN�����3w���� zF)�Y�(ݙb+)�椯AgtF �SU<'I�6u�Y��t����6�'�fU�͊T~T��X��Yu��T�*��M���^x,�%U�0N��،C
����5�����W	D3��/��{�)E�Un�����2�]jE)e6����,������>�rL���z�����v�.�<)����fg0���P��v5�?Ev���pB�u��:$m��Hd�k�/P+?�}�������2�_��f�����w��w��qV"*a!�Xw�9��4��Tt�I�GB��N��3ƻ��1�������z;�L3U�6.0�����?K��~P%�5�w
�% S!��!��AtK2ǘ;��0l�h@H]��E۳��X���yٱ|ĩG�:�.��, ;�RPt��ϙ�zI�h���6���&������I2.�h��2�w��"4Y>�^�l(uńo�殴1?"۩�ߝ��,�"��m��7�C穻�oih8���'� h�J��1����IY� ^�b�UM�d�[�@'ֈ���;���\��7�P�b����.�hmb�NcY�b�<%6��8hL�"I�R� �?����/�����n�P?,I'�+�4\>��������#��!V�6�Vi����p*Sv[=���<؈l�oR�@��ޑ��+!��K!45�C�?`��~ưP��>�����6(��\�
m �UՖ;�