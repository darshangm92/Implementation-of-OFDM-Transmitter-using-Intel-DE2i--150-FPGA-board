��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�������N�4@S�y���zM�|=�ٜ�K㪼"���p�A7W�JIvw߅� �of��Tg}W�t��8�ɺ4َ*��iYJ��$-��m%w'k
auˮ��:��/��ڛ�1�)m;���05�5��>c{
�B&����I� ��@�;�� �R���@g�e�)�Z"�qm��
���ޞ��5+��IB�XeV�M�Y,�ǉ�Z���ꚹ6K�L��*�:7�	X|0��T����$����
�w�q����;4񧃷
�.>r�V#P��<z�-K����A�},�`DUK{��E�ճ�vF�nh}2тM�.@�o�	ȫ�Y�	Y�\x�!v�(�Ρz��#�``ɘ�hڦ����c�f.&���f��]+�uk�� df�[ˈv�<����"�U�=w䭝x�j(���I�������P���V�	2o�%�J���p#���	�X0o��\�IW��ܖ�+}s�Is!H��k`ݠ;R�F���׆;Gug�w��9ˌ/
c�O�EZ�ߑ��@Y�V�c����l�0����\I��y��D��A�iKP8���r����
1���$'�EG��?�~x�Ӷ5�眞���B���L;�~��*m#��8i�}��4�(F_���Էc�ʰ�_�:F��:��cT��q
���;i�Q^��@���ޤ�	�,8� ���0���CGa0�:p��f5{�-�@1  Ȩ��*:���mQ`T�����ȴ3����Ji��G^㓰��<j��P+�N~���.���zJf�y�-��,��iZ�p��.��[ N	��YQ��w�z��-O�꬘��В�������ɵ��`��d�I����O����U/-s������'VZ�'���j�'������	Ē�X���J@i��p����1J�y�)�~G�����^��d�C�Xt����s����m�<�k0nPHl�J߮Y�bR\U2i���(X�����3�4�8��ZWmo�B0.��b����8g��p� -��&۴޿{�� >0y��~}f��Ig�`E�5;��/(��Gu"a���5qc����7�W0V�(�LI���L��yak�W4}�ݩ�vAӰg+�Ǻ�"�^��\p��Q~7 ���,w��s'��rA����� �"Jbn�����{�a��"*1K,���!�v����ˬG�H�⇯�yH!���h,����$������C�f�2�DЯ.�/�#��	�W�����|'Q��jU�pAԆ��N 9�>*�2W�!J�	s�Ŝ����p�럼�a����'���_+�>c�l��<&IR�G�/�`\����5�wS�}�^m�T-�6ߗ�Q;���$�u>je�'<�9�z���E�&��&�^]�L�DF�he���/1&S�O�Fs���^.4+O��E9\0w4V��w�)�}�J�D��PV���J���v��S����	"T�X�U���^Q�N�%ץ�	�nUx4�R����< Nx�X:�[�E#ؑD}��"̓aݎ�[�߿�����('tr�/�/z8)d�j`�N��uT����R��++� �&"u��0x��Ww��-��V��b���B={��dva|��zK�ܬ���O��!�A��H��7�5�O��ć�*JH���!��;���%��{N��� q��}�Bg\H�{%��-�@:$n5YZL��Qk���R�ID�~&�-پM�hin�MѢO-���"#�g�:�r���n�C��5@P��u�q��;�1���N#=xܚ��&}	�]?��]�tD��n��`��D����������;O��[�c�4rD��9q����|��tC��EB�_�_$^֕�V�>���ƣO�ph�m�O���� **����ET!Z��Q�W.�ɍ߲@��{S��0�����K�y�X<dT��?�@n�n����T,���TW^Su[8� �m��&�.�	%�* R�!D��`�Z|ce0�Ï�n���G�\���"|�]�Xτ�!�潸eQ.]����~iX�������Βb�V�,��I��y�W��Y�js��¾�X����C�y��g�ny�MWκ�ӏ���Ji���9�gGM�b�3�@c ٲ�E��0h�걳b�@���X������8|��q^�;ō|"�B<f:��H��,��>��R�ψ<UB��E��O�2u�i�t,*u\��N���Pj�N�/k� �D��ye��|v��`9X6���vArmYK�&2k���A� Z��(�zE���͑d<�@z�s6EtJ_�ý_!��4�����z>���]�\��"��de�B�P�$���V�1}����s簼�4c'��QB^Br���djmۼd]n�1�\�d�ZAu��C���Y۩��U��5��J����*��f��rl����u�<�e�w]�K�$�lf�1���uO&��F�*>��~k��pf����z�����T���)�s5=�����x�#[ΓӰ�BPb���Fϋ��o������=���YJ�������0�����tp����)� ����l~���k0�AmL��\��'��_�1p:��8o�0��PrX�1���L�]U��gH2~J�}�L>��c\�N���$�̪^^��� [<�AD6�8�V=31+n����` $��[?��s�[���������g ����b�j߈U��~k|W��?_�@�J�y���B_���6ϥr�<&��έ2W!S5�� �C��z�aXq��ѱ��W�L���������}���kG� ���q�\�H��6O(q g>+Ȏ�b(R���!o�cYG�j0��jZ�Ⱦ��.�Nzk��gt�iш�q�%}�L�:�2ʘ)�\.�V�zj�B�b�}���r�g$�]*Z����4-�J����D��}�a��b bU6՚���@��Ɉm͵��6@�=NÄx��MO���C��G�zQ��x�=vM��N^X͛��$�Я�U�MeR�Zg"/or�s�{z�z>������#y�c�[ٺİl���_G.��M� �@렘N�U?�r8?������5�E�R��׆�Tڝ����4�8��ޡi�hr9xG08dЌ�/g�r�8<�E}�
Y,��6�OU�p��to�C
pLPG���hƗ�2ʣR�{&�f蒊��e��������n(j>폸`\�Bg"�B��D̊�f,����!��L��s�a:�D=�׌��s��iz�a�r9�};w �;�dc����Göņ=�L�Wk_���;fT��Z���Y�����"�Ȉ�K
�N�JEibpA^P���XA�&>W�����v��� U�&%f�y���v�&��TB���3�<�"��Th?�4i���;��Rj�x��Ur�ugK%�v��ȟH@�M���4/�+��r����	p^�+p�;*.j���I��LPႨ�cF���ǇQ0�H3Ch\9��P��ҠI���'('�� �(l}�ѽz� ��;x�����5�_�d|O��^rXآƉ�=D���(�gOgq�ØbIiCCϪ$�Q�+.c���Cj̃�/z�������"�*6������kun]ٖ��JEH�z��t�������i߱d�� ���LW���αL@��: �U��c�9�Wdm�D4S�zx��W�Sl�|�ъuL��~aV�LG\!+mPY<�m ��L(\};�JF�����*��kۍ~��Hv��$��+�Q6p0��;��� W��L�-��h�t��G�(��"|7tB'U��Q��oq�˘@D2Aɫ���&�uOa��Z����# �b����'��c��� s�8+�-��!2�
��h��F��E9�w�/���\��f5PHl�
є\P�����U0%�z�֫����GP���M��\}�������D�fFѰ@k*���[+\����?����"Bͪ��IU�)
(�l;]��0wnx��̣�#�UY���� _/0�(՝��d�Y"O5�%��,��n�a���7���z��F��Nd�L
=H��#�0qIWb�/�5-����l}��}
*us<d�
. ��l��vG�h����a�����U	�|��u[����5u�f�F�Μ�1�����im��!
t�׊��=���W���s������ե����AeUe?�"�Z�.��}˓627=�?y|p���B�h;�2B��
`.&�gjG��d�D=Ug�e�m�W0�_��4�!?MSn�I���;0��Ԥ���$M�"��g5~�R?�_�#,)L
$^X"� �P�)���CBc�J�Q�ZGt
�fzY�Pc��3����1��Ys'�������;+��<�aA`Ȱ����#�Ѵ=�"��q�Ӓ� =P�Gm>x��5�����{�94���6��8��E�*�P ��ؒ̄��s�����8��ߋ�������1��lTb��Y�u�^4�V���n	�&e緬��N�n��ķ������Y\m�H�`B+�4H�p�;�'��Oŧ������w�|�l��-o��^�:�����HV�0��&�g�b�>�4\kF#��/����f�{����}�E�`�GN'��&���/πn6�Bس�����`Ӛ�W�dy�\�i��\	�#�R����xť��c�R(� �f+;.(#O��;������u�𸭑�~P_$b�I���V"�����P
#�"���^�ꀡ2߶UC`6�8�$�6J������(-ғh�
��\�>���`��Q۩FQ��y٫�G_ޛ
p�/['0� �!��SM�p�����lj֬ǭԚI�/��E��~�Xn�G��^(�\��$�;��!�u>�Z��~��5�P��
l� g�}�X�d�h�����Z�Ac��M�����0���H�s��/Z�tf�!Fw�l51 ���ޤ(�~~vt3���/I�>�܏���ar}w����v��q+H6\�@�9X4/�h�{!~�+�+-�Z���(�y���K���$8��䁜�#�q1Fh�h��
�����@�ɜ��aK��*#c4R�i�SsK��fY���a�ou�0�Wxį��ȫ�;�d��.Ȫb���U`0��b���]�B��̌�2�- #��2�	��m���E��	���c�{x6�JV�l{� ��ڃ|G�*ꠓS��pӇiZ
����Fk"��:E�#b�h�d���9�?����b4�&sv-��4�Q�`[Oyb�G&a��B���B��:Ӛ��c��Śȟ5��ay�"��#5�V��R1���҉T��p�N�(Ȭ��/�	�$�h�&�(�+���C gJ|J�}��d�G96�ޫ~��`?Md���.�]���pe�@D�8G��:!"rK�0�(S���U3�����������Ī��!���ş�K�a������Bk�J��3�KR����"�y5�ZD�as�W��3Kd����фk�,�v�JR:�p�����R�x�IO�(�d�Z?�t�"���}���;V�f�L��!)Ozb21�k p�(h�����P���2ƒ��l�CoV���1���GQ����<Ʉ�oᶞXuD3�@���B�ۊd2�����"{��#��� �G������wAh�����WL�+@&vjn��g8Ho�B�f\���/��.�m�gH�q�e3�<E"լ����I|���B��Vb���/��J�ʈ�,���L�����ug���s����j�ә�l��puk* Jz�F>����lY̡`�= ���^Ϊ@٭k�e��q������	�T���4�STh5ֈt�1�8�j�+Ddl����q� ����t"P���m:]��������"W���a����r��ċ?"j!_dC�G��R�>y�pt[ؒ��w�UR-��U;U�xW���2�qcјֳN�R�̴�3I��Oo�$D��|���^?���#�FĠɴ��
@�1�쐺7tR�J��:�@�0���ڿ逐��C�z[9|���i�\8��$jz�����%��
�?x�Ta��^���<>G0��#�M�x]`����-0�y�!p �� \�����l��NX|�M�0�����V,�=S���]���Dʡu�g͠3�\^�u��l���!�:C�l�+�\9��|l��<490��/R��#JO��]�t�%iNfZ���p��g�>�D��ő��[���z�?m����K"|m�1���À�&�D��ä�����Hm�g����bO;g�a���:1�O澓��Bh���m��R+^��멠�ÿ�7ed/9���b���<��/]�1Ǘ3����d�e(׫tJ�D��A��2σ��r���=����%�E-������H��r>z=2�&������a��o泽XāZF�ݢZ#dB�j����MO3jL��ݓ�J1f`��S����L�e9%X�[�p�T�0g��M�'��+��r|W[��'�p�t���5� XF�s�IW
�R>6ր���h]K�����9�C��9�c�=�T(���0!dG�lh�J�~��:�@(�K�e�N�@��%�8��V��AA�t��AWQ����ՠ���Ee첕��D>Im����C�S6Ů{��}r#�^���_�4�u1��X��q���n�����=�� RT�)�����	M�	��鳸���=2�T���� ���B��a�����ŏ�g{קR;Ob5�v���yQR�*�*�A�>��A7���vI�}����
׊���9>�R�.n��vu�!N��-�R���?*��>P�D���}7c8��Y^�\�4�
��p���tXE��,�b�R�I#D>s9g:�f'IV�_�x�a��� �
T�g@��B��R�<���1�'yC[�]�
s_B�f<���,l,�g�����=����#�33�N��Z���Ÿ^���O�1�G,�����V���1����n����Nd��T�z%#�T��e�d�P��wcP�Wx��A��q������VN?�WL�a�j���bǼ��o��np{:��'���p3�l�*�׭7F$�<�,H�%s�-�u}��qfp���KI9��	��	�DOQ���b=3�^�֎>'��M�����8B���OӬL����n�N��;ι����"�ۤ'�� ����u�y�i�2�9bS�|8Y[�F���|H[9�X�{G�&���0� �8_�1t
�!k��D�[~��k	U��W�߂�����:���@Ts˻�i:����f��[�w�M����.�;'��+��=\��X:$Ӷ��������`����މ��������Z�V4}�G��w��~w|�I2��P�@3���
5"���$�	�7]��a;h���+�ؤ5�b���̸�L�8P� �t�-g ��]���=7�����,����!�$���� �LS��t���_4�ge�~�3c�r������B��l������]E�b�.������½[��֏S�I�\��"�qc��~�;�k*�-��6CBτ�@���~l,6e�ǀbڼ���*�*sC�}�)����A�Uk��u�Wr��	��q��p}B�͘f�O��jR��h�g �����7���W7X�9�u�d�ƐI LԉW��R5�,�u^�]�b×S�-[�q:?;/����V��o��
RO0��3q�<}�!�Б7}��m�p�9�#Q�c� ����{lA�������~s5ز�5�����ګ٢��J �{���F2#b�ͨx��&�𳇳hⱛ��g���"[�����h������78����f"ҾqΏc�':������0-�n®���N�ti���4i�4sl�����ص޹�A����"�<�^1���SZ?g��*����O�/d�%�ɶ�w@�=y��p��8�%|�(w�nJ�7�w'�U�� ���w�1)ڼ 0���� e܈�7����e�c��T��iQ��8��%ק �ցg�V��b��s�vHm+�ƙ_���|h:k*�~²M��y��A����A��v����?��<5Y\���d E��)''~zr?$ۂ=�I+�����b Z�=ԃb2ư�OY��� s���oy�0��7��*�è�61H3Tod�#�/�*�ʬzRHF:{�N1H��\�8�&xػ�W�H�ގ����[�¼mD���y��Hu�����li�g�)��6�"  ���v��X9o�j~�rq=��a��D�����nyXv!'��m��X'8�-��K�d�"��Օ�&����Z�cj��˛�Dl���%3���8�w#QpĚ����W�~��f5�ڵœE���`m&�$��o�-1Nj����ֵ!��@��u
\���8!4�ņ��%s�&��36�<.sNOA����bC�oI)v<���0M��T��#N�<ʻP�s�ſљ�C+3�"��"����3���AL��A&;�铑J b'J$���)Fz�0����!f�X���9�^�6尩�x���k�����֗�73E�䱚�� N,��BL f7F.-��Vh��Ѽ�f��9�����m��C̈��D C?��",�#���%3R������h������+��d���(A^	m���1�����,m�	|�EY�;�כ;���5�Ȥ�T�<"�a-�e6�BY�Y@͒��ýꅥ�ey�(�z�
��a_��w�t�Y��	���f�\��>W�>~m��Y�[���7p4�:�L3�s�#��������C��!'�j|.�߀U��$H�[ǎk9^��5f�ۻ��'BhZ�lO�������+�pz�t.��_����F�A��(	!/XU�+�<T!�Pà*���K�T(�t�Ͱ���K����S�y��ܖ�ק�+R*���H�1Jƥ��0	d1f�eG��I
��1��10�t�2��6Ѝ�1�{��4��>}Ȇ�D� Z�j.�A�G�{� 9�����F,&�{ؓ�Ia���f��y�{x��Є��b��5�������8ۻ����#O���P��f,�o�����8&��U����]�b6~/�W���"����6;9ݙ�V��e��NW3c�R�$��I$�`���s˯5Ŋ��R�xaq�l���qKi��;#Ӳb��
�yv�l�	%�xVv�(�W��޵���Y��W��RV����y���u�W��Mɸ�v�>Uq��.J�>��[|	�T�@����F��PQ�.h�{�ۺ�����HN�J�5�P��jx�|�PW���;��܁:,��{��@��TB�����:\��L a�t����u���@+ς(�_�|��K��t�[�u𕸽؈Q�k�����
�����M�w�j���9������
���o՗'Ln.v�Z�Q�TJ�b̭˱�HG����py>-�P�u}1Ƿ'n�ùR��}�q����E�:ș�� ���4�$-ô�@X'�a�Cv`D��`����"m���/�zѤ)�Q�Q��˨��q�Af3JM�V�����i��w�����,qOv�#6B�+-$��P���"����|�E�3ֶ	���Ih�ҀD\��[�;�H��@9A'��Y5���p��H~����X����ͭ�Bqi�.��q�������4�]�֥��H�Ʒɟ�ىx���X�z�P���0�(m�?���8��}F�c���Q�3��.�R�F�n������j�%����5J\x�{$�6-�gdk֌��9�����#�4'ˇoS} |iƵ9���:8�X��E|�*�=2>���Ȇ�'8��=D�AX��z|]��s)΂Y��N'��C�]��L:�@�mJ������]Wl.�2_@2�Dg�(�u­-��*��kb����f�2s%#�ys����n�
�
P{���M����톌Mf�@�Zo��TE"��}`8L�"�)�it�
��tB|	�˳5�Q�1���:�2�;`�:<qc��t�m�S��
��V}��24���˽�O��;�7��d	��Ό����`Kv�UP��.$�m�l8	#l�<��D^�s���ª�}����j��D��V�Ή���#�L']�'�f�wJ�Կ҈��_�+�u{�\JB�Su�:e��'E�������gXDP�7�<'Zmׅ*�����	�d� �=k����&��=���4� ����r8u��!�z��������+��zsA(ɼ� h �+�BրUP������-�/�9>�˄�FO0v�ÞKz���P/����Aص%�콍�v�w3ʾ\�#0�eV�� (��+z��JHl�����$\w�v��	{뼓5�?�g���1��9~ͦ��v0���i�@?A��ŇgN <wﯜ�i�W��&,u��v�Z�z���H�68w*��/Nα���X?�jf̵��O�Qsk���قM�֍�� ��yEsb=i��N:��+�%��
zsxJ��r���� %X������A*�z)����.�Gﰱ�˛�$O����Q�+�2��4�0�W����P��i�'	^�,��8b*��k�, y
Hd�-���o���,���6���kGм�r7+A����g�_@����Żx�i>�H��� P�>c�˯4@g��塶S�������3ڢ�]���q�U��:��mЪ���j��S�[�NF��(jt�'E���,Q�CA�x�.qjA�ԓ�"n'��;eŗ��Ju�I��;"p-Y�;*,��":P�����/E����0���c�J޽<�n?6="PK�4MƟ�N�C�0ٲe�4!HV����0�fQ��Eǭ�:�����*����C9���>�i�=��H�h:��T�HQ���ԏT�L�25M"�<;� X�l���ɼ-����0�Xis���Hv1qtT>�k�4�M�>�x�g���md������Wf%B^f9��xY8��pg�J��+�ɋ8C@�S��$R�E�2���R*H�l6��P�p}'x!�8��V襁s���f)t��G�I�7��֊��E��*��i�gj��T�+�sԘ��|�L���JB���Foy̓�2߲�qW�g�ٵ4^�J����w����?;YY�g�LsG%���}Bt��7���?�C��攤/|�jy z��2��k��/� �؞/��ӑ��z7	[���rͭ���~C&�h��6e-/��/��A}���Yp�c�O"ۙc��T��3˅�:���s����/2�z��I���ހơ��EA^%�����Sr�K2�Q��c��	
M	b 7�x�81Z�|����� ���}������ؑ�Ѽ��i��i�ǋQ�&�Nkس�d�H�������0	���?�����P���o+4��]\�g�@�?�ď��Qb26u�'�n��P+m����U�4~hֱDNږC!b4��Rs�����Jє\^ �m/坠����/㸗�[C���!���ȠsB:
_�	�������Jn��<U�e}�Y1��V�Ҭ>���z"�u;�֖"N/�	R���N�N��8�<��x��^N�(v�#�/ h��I�C*�qk���F7H�b/�S��
lNć{�n� ʵȕ%���Pb_��n{�ٯN�& u_����&��}������;�
��gs7�xx���/s������Jw<w��PྎXi���i�a�ѡ���$b~�8s��r=����h/��v7S�]%*��^�2� PLF3��7��^y'8'm���u�vR(�uh��ж�QL`���Z�=����uaY{�K��ۘ1�M9��q����T����v屏�H��z�C ���O!���2�I�+̀F>�W�&����󾄆���{F4�10y�Ht�=���XI`57⣡����F� �0���EieE@��Ȅ6,�9�t��9ϔ��@��r�Tk�f�e��T�o%�-��m|�%X��(��jT/�R�E��r����	�>���vS�Yȫv:=ڙ#}��8�0	��R�1�����ܨ��&�g��m�~:v���#?��4�#b�h\tkIݘ�:c�)�u�a�h��������RiIn`�Ҁ�Iᱼ�]��i�����#��x@���b(�.��9[5xC���v�=
7�뎍\s���m^Cy��{��)]D��t0w�B�H���^�?^����������7,q��q��4��b�P4��L�%����Ec����@E1� !��x�@*��;�U�&1�1)xu�\������ 
U�I6�mtW��z@��!'��uΧ+���\��$��+��;��x~iPNz�b��ꬖtkw��f|j�]=d�����>�����EH�J�s��V>�3����h����p�^��ɩ�f����D��?*���(���_!���g�2�MX�o?{Q���e z��3��U��O�b�
I��V�M���ç�
꽕����Fy�S���TSȩY�ËtH���e>��K�zeg�x����#6CJF̒n��!x~�`�
�ң����8�4 G�}��)�]Ly{�^n�%|�3^E�~N����0�M�H;+�7<��`���3��U��AQ�j8s����	`q��7Da&6m�#(m5Xj~����y*���Wy���~8F�ТÝ�$���&��DP#�Ж�xC�#��G��S�Z8l���p�Ň��r��; "�w��h:��*�1N˜��W\jJ!B�'613�f<�T|�ȧü�m�#���V-p������_BŔ����0����ˌ���o��K���j\�_;�A�&�E@<�ΒZ�) ��l2�}:��4ǒ��v���?\�E��4:�K�7*g��ؠ��v<'
�J>���a�<#�����
VO���kDǦ��W�$�I�2jK��Dp���%Dխe�\�?��M� Y L�Z0�Yw����ؗ���J�M.w_�cͩ����n��Y�u��T�&G�96��;��s'��XcE�LҹQ�N��pb�@W2�>f!煛_@�W�֓����NI�#ʱa�P��|����T�'>ۼNs��ͲK�A ����TaڥSV;?x�$&��D��fId�e��U�1�~�r�Q0JSb��ó�H���O� �҂��G��V�18[��C�Ȋ�������{�L8��l\i������<�����/� �XASDim}1��������u����)��)��O�:w"��Ea �����J-p�����D�fۘc�sּ�t�L�K���V�'Hd��t�����{���G;�fԎ��F8�h(cUq�bc�Z4����7�_��ïjq77+�j��d����K�.�q��f�c�PK���9�K��v^���{,��X+��<�z�)��F RSK�q���x7��?��&P�8��2M��|3f����	�h�wo)"���eS��i��R��y I4>e�u�`�?7+�Y����*�y�46�#��n�3�d9��(�3���Vhe7��<�ݏ ��U�|AE�wL�?�爾��g�e����d�]��kI�}f~�U���'�t�/��*$��|C��5PO�����#!8W�Up��+�,P%my|w���+o�V`�ȳ�e.�8�Y�x����1��T�&�bǚӓm� ��M���;�bnm�#��L�8c�g	��8��8WI'I	2��b�bT�Xaף�m�TM��`-����fFF��R�TOf[�ǽq���Q��+�-*��[�݌jd��ȕ�v�V�"�L�Q�Mc���<'; z�C�� \J��!�7�۹c��	�pm�H&�:c�`�#hd��j��Z�F��� ,��X��������;�gj\/�_Z��T~��`�4ې[�儯�5;�||����*!�#<���Y�(�8��V���a�j�щc��ނY��2ဍ�:UnCPV[�9�Go��a����.?����C�\Q�d�Q5x|�cE���:κ1Ҵ�ɫ9
�"����S8��>q���@Hy����q�+�SJ�|Nv��.��QlʺI�I*܄�q�$"{��4:�.3	��<��s%����&�tc �O�}���g�3���ڢ=p���Ҡ}h������u^����貓6���5>���^x�d��  ���]Oh@X�J���lM�$k�w��GZ���<|&����E���Ʒ �f��8�PR�ˑeW�������1����ɝ�!]��\:]���hc�M�h�E�y�MBܑ�!����X�����x-��뤟��G�����2��M'7��P�T��{�ky������6�'��ғ��k�#�<��Y+ ;��-��`T�o����,��Ρ\���6,���?��y��@#�Ӷ�
��G�(	��60VU��!�6q]�Ƨ�T����]���ݞ��q
�o�	*�hz�Ȯ�b>��4�Ln���;��܈��X[NBq���*�� �#�	�mQ�`��WύN�EWl[_�ׂ�ٯ��l>~3�u�}��/����j�"�����uRӚ��X&۹
�a�rS[˥��L��m�څ��	�^L�f����Y�B�؎[�P�~~IL��9yNf��XCY��P���pW�s�t�Q�E�F�PxD��8�4��6܏�L�W:�~}1xR"��y+B��;,MN����JgB�E���&��.���Y����������n3�p�l�'$��i�bI�,�PG\���.U��huYU�gwS��!��(�@����1=W��ӲM+����f^��A���x	��eօ�-���`H\����Պ�/��`��N�E�m�z������y�o�]f+�nZ+�S��Ș�=aZ9���(4�^ɶi���Ηct�&wX' ��)��w�$L�l��R:�ӞnxY�>�zj���C�����o$W�ǀ�C�xoN�"��E�A�=�J�JȟW���?*����r�ëX���T�]'IF��e����?���-����f�`/���$��NK��m��veL��/=!k��R@ޝX�dw�ވ&���(MB~��\Ϫ��0���A�H��VÚt�5o/$Г�x"�h��[�2K�C�>a���b�"� *C.�	�L�Hg~�ϔ���3�-�N�O5�k��¤ �D��>�@YJ�+%� >c�/�Q�~+={U(ǩ}tzt�Uv�F�>������j�V۱���
� ?亂�V�S�G+�ι��] �[q�Kr|�-^�&k���*%�`��#��⧀��`�؀��P�˱8��Q�9k6%r[��D�m��3�H0Y���ș�5p��١��RV�k�1�+�O%3��"C���ǟ_v���v���v|	�)j��{\�9u��Vo�q�k𞟄;��b4���z^~=��)�-���&���KmDG=):o�:�H�@m����f������Y�Q&3eխ� ��~ =���O5� ���swm�e�R�/o�m�P�k�`k����o�@ ��L���(>�\�����A�Dm�6�������7�"6�.t!�	�v���]Z����IU�ѬI��V9Gp��hb��D.�/3�h����5�^n�����n�m(2�r�
��f��c:lǒ�m�ք�����^��3,GS;��j˨��v_~��Y�-�ﮆ�����;����#=Mt)x�a���U%���� � �Q��K,նGl�T<���S�X�	�%C�-���]]��VM�f�L���%�����4w�j�[�ɴ�/�Bʂ�N,��ԃ�^g�<�)ߜ$\�8�]��W]Fsٷ?�*_��y��fe�'ʽD�o��������P-]�����%�퇸�ۀy�e�H�R!܄�G%\��>��y��9	�S���Π4�<�s�.%k}���8�������!Ѳ�s�qw;�,�$$�h+�8M���1v�M�(�I��A� b���SV7��D�*�����.A�Z�Ëc�˽�>7W���p�qQ�~�uz�5_�מ(�_��G�'-��1A�1��S=�U��yOü�^�Q���٭;��fF7cY�����'�ef\VM&}�h���U�+yA�+�v�Mp����%[c<��/t^�`	����yj47W�����Z�x,<���M^��U����a�!&8Y%�Ƚ� ��\/TN�Jq�^�-��1��*�SA�^\[�1)L�i�Gb(�Q�I���<�$�Bũ=��ɵ��q[e��r�~���V�77+Pw�䞃Ǡ� tt.eh�2��*¹�祐n!-p��Ayr�@4��r��^@ǋ�婭ʈ9?
�њ���Xj���r��0��D	�1k�O� L)��ҳ>�?�Rr��*��Zx��E����(��ϝ�\���Ε���lćݡۅ'����R�n4��'8X�߁�V������t�H�#��
a�B�*1�` �8p�Gk������:����ĬĨ�{�V����������گ���ى+�R:�v��Bd�o����ɶ?l}2��4����,�坯�A�k���bQq�"MC��ד.�aYilw�A�����O��"
8#���c!D;#a;tg�h��D�*z�՝�b���IH=�m-5�'b1B,�n��@N]��!��Z� �H����j��ͺ�Iz���	h�T�ֆ��K�h����]�-��&�|��l8�Ďt�v=��M�ynP�v����63Qz7��W����"����$���%�y���\����;	�ߢ�姧�JN<���T������F��D4�f�Q��
��rnT�b��I9J�ݝ�E?�"nq�����6��FoX��xA��������+��!���y�[�5�+!X${Uo;K��v1�͔��Z|
�������-Rd��8�$�e�w2��?׭�w6jn4^�A��/��M�z�b�Է:����S�*�ݣTydyؚ�B�^�Y?�x!�Sn�i+Sz�)+`���6�������Э(ho?-`9+L�l�e��\V<��q|'Dz�_�|����z`6`?j<��J�/o�-t�Q�n!����*����7�fB#E�:��MD`lK<�|Y�ϫ��΋�u9��Z)�ſ��g��V�T��I�5M����y�2?1���w�
�	'�4c�����]� +��ɌB�<̯�W���1��@�`W��9�R�U&i�F��9��C1��c�4lN�&:Q��jG�~���>D��j��Ŧ�fXX�
�N��)�?�_�M10�E؇'c��Ά��F~��F��L/�~������ￎ��}k#��<�FM�x3�O���V���ʣ ցd���f�(*����SCǶ�,�ӵL�'��w��?]����^��᜝��bŚ	����:6ˍvŰ�g�G��Zj<�6�C!���.sꈘ�*,H��$�v�D�y�-"�ϵ����$v���t��Q��4ʹ�0X�#l�ɑ�nÄ3�q�%/�]�
�,>�r�`?��h%)G����0�����TjO!���6��#E�
!<b��7���@`�C_����e�܉��:k�`|7�(e8�S�@����!"��(QO����#����U�nm�zx��-&�4
*���7N����E:Qk(�W�8"��>��Kd4$�w��ÿ��w��F�?�Zvk����A�6��'�J*ʣo�eC���'��6�	���a�m���YQUS�P0�4б)��GuB��M;Q�C��Q���V.�C�9��ܮIT���V.c�Q`�*��"�\2u��by�'�&&�N�������������v�^[>��	�X4Ҭ>^�iG��1���Ww�~��\����_�
��P�)_Oמ����dz^T~>���7%9�
LS�i��@:���I(��ڭ@A�h�{U}��*�y���6��N��ҠF��&�-A}��XRd>|7fUK��qɉ5��0��U(jX;�B[�>H�Ҿ���\���8˅_��Pm�쳬�@���O�-z[�7_T7�P�톭�d���Ӆ[�g��#6����w��R���WL�5
���e0���W��L>�~�j��V�jٌM���'9b��1��BI���M�P�!2���{�#������5h�ގ)b�_�����"��Y�8g�� ��% s�><_��~ ��l���6�0 �C2�{p/�����D�]�48�'�\�����Aa���	���W�Q�ua�sCB��~ݿ��G�u�b�Ч����9i؊c��[��^��C���	�Ĺ9�A�]�&��?@�W~Q�@
s7;4��s���;�j��3�����v�c˿�mFMF9'�g����_u�^�����s��;���b�Q�3�{���?o�Í�_���HM��'�Q�7�թ �:���Ϸ�����!<�p�<�S�n�9%�ҩ/('���t6�p�:̵�W��5��Gf��f5D�_����%����F�����[��<J���`UӋ:��.����//@"��{`pՖ��ף��,1Ѡ�#QҼr7˿i��@��y!G���9��i��7��U����]n������'��Z
���V��������}�ڿ�m�����G~Lj�&���Ԭ��a89%X�N��1>Yh��T�7�٣k�[�x���~/�`��]]uSt�گ�|��rjFl��o�F��^6D��1��8i��6O��8]3�_k���j+W|e��)I�U�s �G���PYDw�=UlZ���d�cT�ړ��4�,�QE��44I�%ur��[�` �x�J=/����<�?I�*3�)	� �tF{�]�Iy����o[#á�ʏ��c�_bXQs�1ж��G���C�6mM��T�VǏ���u�Lÿ:����^�Z��r��*���>���T�|W��(���5���.����X�5�+)��.�2�u�Kd�Ȗ9:#�i����c�c��e��d����εg;�@�����:-���YxGd�o�F�psur���?3̂�`�w��c�����.�ZuA��(���)̩��ھD�\LM�>D*��@��T��ސ-A~��t"�˚!�*�K(�䮻���a}&�Ru������!��h:����=���[���ۊ	�7��6���H F��89�8�-�=s�����F�]4��t�5������^ˤlwҕƟ��;$��m5O�Nvt���l��G𢚩+++#�'���"v��g��z}��	QF\Ne�ѷ��&��� P#����a�㛱#|ˆ��{�����M	��~µ0��k�V	������*�>}���cY���x8E�ئێ|e�j�H�g`1�*b�>TQj�|�ِ�@!�(:o�G���*OEE��G|C�����8�k�W����6�u�I I5����\,S�Iw�QZ�0LDԶ�,�}��1:�f(Otd +}ݶ��Ƚu�m/8��8��;��}�.����T�h��}rM��Ƌw��d�
�l%V[jw�ނ
nk�%��d��.�Mt��Z��9�N��������eGWF=\j,�,f�=�H:$hy�YV�N-�Ϯ+�ɝš�����l���\)�^ɾaF�'��L`���5����\�z��_�9JL�>�/U�@�b�ȕTYc�|(;�\����L��ь�#�,X���+��4*q��E}����8m����{"!���s�{�If�q駐�M|����T	���7(���6�y̭^�V�G�Y�2�d^�6~����:����
<����#�]*����8�<�^#�Z�>A ���J
�/HzY�w��锋t�EM��=@���͙��U���>�mH����Ř2�Pa��M$��.�H�9D!����[z��`C����ތ��o�=��G5�r0�똳�D���:s�w���Lv=mxz4Z��N�$W<�c>��P=ߡ�v�[̴���@6YI����﷌/Dׁ�~�m����-�����a�2�>��5����:����yX0-㵇]�&�^ѲnW�᯼���A=�銣S�G��`��FVy�q�_��O��mܳ�xVWXVw��=a��gQ��>��b��?�bI\�X��]��]�����W?*�f�F�
n���2'�I� YMc�O��T���M�����'J����%Q�ԴSU`e|�q���䦨�?k�v�kA<[T�*�_5�@�J�@���|u_;�B�L�i����1���D���C�ic�%�� *b�*��F/	���4`��m�C�s,h�x2��\�&% %�OK�Z��.�L���f��k�?ו� ����t/�@X���*��#)Am�;E�s⼲�)ӄq&���fsl78G�:���\�p�l���tR�Ďϕ�5�XbQr��j#�!8[)�z���/���c���P��\���p�[��y^��� v^����0O�����?1�'�Z��Ê����h�=���{�	�/6Ӫ��iu�B~zzOC|ϑ�(�K��t��Լ�T�O�U�J��ͽ7�ع:4L����^|[XX�S�jQ�f��+U��J��ŽbV���ڜFv��n�K�u��i)��*�����P@f�m������!��+�gnf����7G3���Y{�:��	L��F�U%���j��l������DhS��f�+ΕE��^ρ�PW��'")0���a���P�&�.�<<�߁78Ј���{�+�.�)Zi��-�����$���D�*� ����	.�'-I����'����b����s"�8���U�DZ�p"qnL��! �PH�6F�/̰�<^���Sf`L_7���i&h�)<�����Q�$�o��6��������K��\�ժ�2���Lʜ��b�x�k��R��%��x���$���K�'���V$5��H�����hW?VG	��7�4���>@o�ܰǼ?/��&��;}Ϯ��ʱZ���oɘ훙�v��}��Bn`&�,����0Y��zHXmfw(`A�� X����k��(�aL��\J*Bj0��F7"�� @F��ǎ�E��ɮ�R��<��'"��2���YѾq�ǭG� �Kc�5 �_7��jbx~��[�bR	�qN}zz+6�"xI�����|����ֻb���w�vX��7�,?�P	N�����Lr&�LK$�.k4�J��������C���h/ ��嘬FC��_�ez4�o�{�WsRo��s��i^�M�(��ߢ�Ed�$^R(��ex鎈�A��IDIh,����v1�����ލ�Z���ʯ|R��D6�d�����N�x��>��b&�M_���I��;f�<�{���*vآ���\e��xF�s��B0�4��YY���P�W!��֖P�V_OR9������f7��|=)"���>fX^�}S#!� d������9�.�Օ��o��V��yd�Ӭ;��ߗ�L@��/w�N�!}����Ő���o��+0��L�Ҏ�+�a�B0qV0 y'����K�ʁ��]}�Q�#&#�{R����$��G�:��`�T%�4�NR����ך8W�sv�Z����m�|��߆��Rv+� ���A�H��5� ���7����]��z\�f�v'���J	��;W��MR�Vo�<U�G<'�_\I3to����El?ǿo�I��F�U�����O}�s�7��	Y1d��&�����Mt��݈s��].��$7|��2��#o��.���ý���!Ԇ!�[����/���P�A��JUm���<���G�����Bݘ�X����I~��lh<�o<���id�
���1
����^�ޕc�bQ�0����XoH��\�)��%Խ�ˁ2+���߸ ���89[��0��K�>2fC�*��ltP��I����Z������_I	7U���-��3�Ca�Ub��l� 	�_�OBv7*R->+3C�&�iV"��Ԁ�,�&�'��A���I�y��x ���μv&	\I�~� y�����C�&sO貲`��3�D�A�L��Ș�<�ߤBYR>�o�zz�3�6r�魪O$�?��CO��I��^ǭ��/�;یR �Rmw�u��O��>Q�ٚKb��Z%�i��<� P<W��Aҽ½�+���IXb
Á��ʯj���  �`��i����x�
O�F֤=���?�ʉW�-2^���1KCSG��0SJ��raT�
�i��x��~Av��b��`�W�M*�>�N��R��ט{�'u�߱Q��V[��uC�����?�?�T�{�>�NA�YU6�{����ԍ(����%{�ͅߔ@qo���,�P��6Vü�n°�u7(���v���y��"h:x��#��e� @������0�����B�<�(�SM��ef<�M�o�:m+j.�29��b;���<�������ܤ�O����@���J��sM7�	[���rW8��8���>{SA+l'�ěw��5��×'���{~�/���8�-�Sf52�.|S�O�hQ�bn���Y�V�_jN?	�'{�k�"��o�M�'R�l��Z.U��0���+SQm@���{=fڧ����㬊����J�9��D����R^@����X"��]�㈎-�n�G���g���=*.[w%#gq5� v�uz��yBB\ʒ;���9�g��_#��.���j���^(��4��:��<���B�@� ��{yaΔ������MϊLؼQps�A �j�2?~ẇt�{��b��޿�K���z���'�f�ĉ����-
V�4�̛���u4E�����&�\MW��~�����T�*ս%DX҇��{
t`)�?)3T������X�~?�"���%q��:�{~����� �%��t$��`�,��~W�#t���� } gj_�������`غ�)�q{�IG���B�&�m߀bl��К�t�Qv�? ��8G�`9q@�j�f��_2�k��\�cJ����VQ���[be�W8����O@�q��N��u-�a���~�h� �7�����!:���NP�櫓/�\*V���va�����ڃ9F��HPxa�%u���ѥV���*���:�3B�������SعA��$�@OF���H +�\�$_�5�yl�Òl�8���#�pd�+�F�f��ܟĦ���F˯P�) Rvd��T�������H�vb��8���G���}Q��Hք�$�=#];J�Y�zx��y����Ҡ�