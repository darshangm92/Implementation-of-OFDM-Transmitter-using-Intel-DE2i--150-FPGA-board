��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����)e���0��q�=� �%e����j�I��4m��b�����u$���r�}s|Ά���EF:�t��c<���n���b}e���p�xn�����V �`��H>��L�F|�җ+x�࠳j�A�I����P�>_T��i���]ޔD�_�l�#��}��R,���>3���&�[����@�J����OA�v���_�츆R��]��+�S,���p�Ю�J�&+�����\Z�Y��}��n����� �Z��}ϮO�'*�,9��^����r5a,��-�&�1�����m%�>��/t?�e���Kz�B�J`	z2l���^���e3�0�9�xc��^\� �T�@�m�*b��y�VI���ڲC�jCi�p3�
�Ʋ����9̸s\��q�oD�
��>�����~�������
@��h�U�&���c	.��<���n!kg�<F��v�+Qd�zrE� Cv�y·݉��cl����Q0�p��.�9��6[��Ƭ:�����i]�l�1"x͓�g��D6�UO�lz�y�B���\�~�>O�Ѯ�`^�a
�Gj���ج��;�I�80�;�~9�#���������V�#:	����b�*�.d� ?�1�W�i0�؇��_V�_FC��*���sD��X��妤���͋?��'����u[ȗ����F:�Yd/�8f�F�Ai#p�f0��W�!|[�:b�0� �����f���������
���h����1;A�?8�{5� �DfJ^�@����-��E˘�<n�h2X�kg*��* ̀۾`�)�M9e;A��p�Vkk"��U+�;C<E}T���m��p(�;-Sm�2�RY�s��c
�M�"/�н�����oHϳ�9R�{<N��Պ"z�*�Dx�n|k��2�6��J��k����Z�Y��Ac�%c������;P@,�5�C(�G]�p�L��|q�:�E��J�I������j3;i�.ݜ5���պ}���L�:�Z�>WP����վ�����ō`�;�u�)`:������BV�A�̻O"O��_=0p4���$�+X���5rC�O�#$D	��k_���0�kw���0�	�@��Kr�Ry���}O��S���F�o�'k��pMa���R
����Eʿ��3���Cr���1��V��/�z���(D{����/nvX�����2��4g��P��⣱���(��fauьR���2�U����@艢��V��1�~�K�x��2缥���~ݧ(A���#Z��P��?(l��dbW��<*���I_���5�V����L0J�E�������K��O�����J�i�!��X��oz���P*�?)Y2&'��M-�(��i��q `�Y��0:�o�8�u��t�٢��#�X-1��*(�~�Ha6��"X����XDӇ���?���ƈ�r�6]���Rӹp�K�!� c+��{핺;.����Q`n_�ֹ�\�
���*~�v��GQ�]q��{ p�H=G�	;����������T|�4)��@�؁�"@�9��j%�>q5��> &��D�m�h򔧍	U/�h�k��\�zpC>��!K]++� 59���QF��\�?/`�ӹ��ۿ+V�sD��E�"��\�ް��(iY�m�
!h2gy��%W�	L�����v6q���8q���{��^߫<�E�DE�7H�8_����$��j�1����c��C��
=FC�daP�^���b5��Θ�-b��'ˣ�By��D�H����/�B�f�*=�J���(Q,ч g��ر;4 ����?}|�s�  f�<� rE2���e
�
#��&�GFVr;���������$%�Г,ꉓ��uL��`���{T�,�
/�S�-�~8N+9;�!Q3����cħ�19��i�ŬFC����f;�;8[�F�]GL�|�Jf
��o��c��I3���UK�Z��rV��I��?�����a�?��c�:K8=�����KH���wω�q��:c�#��N���Q��s1|V����v'�7[3�0��6��uw@I��g=�޷y}�Bͩ�zfU�֊�R77��\m��.ݺ�3�`��N7�����+0mg�
2E��u���&D*6��m�k�����MU��ġ�����E D���Qk���g-&��N��m �,/��wA�	C�4���sQ�@&D^2�r��Ϫ͊�<���2'\�~�'S����5Q쓙�F��1��Da쏁K=�}�v��)���S�<�����|Y�&"�x�Y7ǰs��NUl����C�^� z4�#T>[�9���u���d�ɗK ڥ꫷�����j%p�&� ��^zk�6�ރ�Q���T8�7���Ӏ�=���>�
B�q�=f\.�$�$wGj	D��eI�N!��I� �%M Q��(�wc�'�'Fpա�PϬi�v��gwr�;a1�7��$
�l���@���t���X<(I*ͮ�2n�
� �֕_6��I���
�«R�'Ŋ=�?!��[�:��=?hK���Wh1�\S��Tl���Ka?�D��$�6q�6J��|�&�x9Ą!�B��F��4�u`��F�tQ�Hk�y��k�s�l��ox�x�f#�m�Tj���G�V�}f��k�*o�*izE�K@O��P�����l_�؄�#*f��%<>a��LI{�9�FT}�as�?�u��xFB�
�.�����5�e�J-������=�ĥ	^��A�A�\�yUEhJ�6�L�����;�-��N�A��#z*�������mPp�����7������[#�~�_k���2��>�P��n����RJ����]6]2Z�pd�ɻ�F8�2���d[�hV�u�Dg�ϒ��)ǜ����9�ec��ڈZ�/�T�Iĕk���V�F.�4#��� ��N~��hs#3 ��([�vG�<Q2E:]��{���_#X��P����nǂ<�(L%�o9�41�٭;�j�Yw��a`q�RH�3W���S����n���s_��ݛ�xX�ဆ�����)&���� ���ֻ5��g��_��E[��kQdg���S+�<�Ɯ��܇�&!���}.��B�dه�Yu^ӿ_�r����և#�;D��N��!����]�X�6�t���SV6#*p�\�'�U	#Mmu��~s�G���A*�?&B��L�x�%I9E�!�z�M'^�eҗc�� :��G�+����߳+�'��ʔp �r�����;�G��3ܬQ9[���������X}��?9�\TY���_����پ�`��̈́)��a"����I��
�G:�M��V���C��1����i�	�1�SiϐI,��;��R���d�y��L�F*��W����l�õk�b��H��'����M�����NF ؃#*��׺F��"-��c໒��kkD�����{��V8�A2�_��)��C� L|
d�*HX�xԲj��eS�~�R��1�!y��Q{�e��-��(�f�t1O�G>��N���V��yOg&މR<l8n��O�l�H�U֑�5O��@�m�/
��-P@�<�&�%(����*�m¬�-����tTPVN[!;:��Q��x31񌜔;l�F���T�Ĉ��/��9 *Py��kO<�>�T������uf�H�Rsz�e4�1QأʺN�y,uH��F�V�l��A�vՁk��L�ڱEY��=�s��v'�X멑�wõ+� �L���Ӽ��R��p$���|[W>8�`�z�ˠ�Vb,r"r�xRy�2�1��s��K2�s+p��qX��$s7��/�D��~���1op�v dbbZ����a�}Y�{	�j��>Ҷ���Sc�>�P��:9�N�X���~I��������}�͘?�6��$|���ߚ����79��&�FiFJ#z�L�Ó�Q�1em�v4Q%?!�1���$,�t��FSd/B��LY���!���GC��4���<m�[��Δh7TȆ6���3��{�Y��62Z��cIEI�<�so���$�o�
��SĒi��¼6r�HZont�]_Є�'8�Y\���Q{FrU��O�{���g@nq�r�G*.hZ�w�c-���z�^]����#�w|�5����.��/����6���FqV;��_����Lh�[����ڱb�ػb(u:gGG<��A��n��	���_��;)�W!��q�b�lp��0,�'Ѓ�3\�P`���+nތ2���m��7l����_�@�����������"DƋ�t3+����+�IKҙ������v�J���h�]�z��I�t�h�.hӼ~;�0�ݔ:�-ޖr~�\)��	d����~a���z,��Q&G����1G� ~Nǁ��uF�����0����c	��Nb�-&�\��	���R�~���=�{�M������H�Z��@v	FZ{�:��n��A������L�����+û$A�v2�9-f'�6N���ӐW�T�S�6�c{��Y���C���(�C B����'7�FO:-U��~��jy������?�c $츆16������\�%^���T����7���7�G���V���#�U������S�}�fO�D�WB瘇�䁾6��1�#v�98�|f�ş�#En�p=�B���g�j��_��+�[�)��[�k \�d����E�����e��mZ�
۱"԰j�U��K�-���� ��#k�:B�j����Νrp�Ĵ��q�8��}��������{W(���Q����!	������P�$>-u��s����B{�x��� -��r�e�
�g�s ޞ�Ϯ�����������$/w��A ��<(�):��?93$I��P����'���x��&{��?ZO.�'4ȋ�u���_�s_��2 �; �qR"�#|N��c����+�_�'w�2�D�┎(���L�#:.��"���؜���1Qkϩ~m�}�\6�(t�(4�v�d��l��?��Y�O��,�S�\���wbg���;6�rlG��,wgIJ�}	�(��o{��E3�ҖZ�;2��7 H���gX[RE	���ְ�w�e+�P����ažFM�݈�B(���z;c�ӛ�m|5�My�Cd�����0��}��|�����b�.a�ӣ�?�l��2^r))H�W,L4YQ��<����bw,�q�[M��C��ٹM�n��O�RL�l�X�i���E���3�}N��&ݶ�ӊ��B��L N��<�Pz��+���Ւqq�-R7����	w�'A�V�Uw���$�!�|{�p�E���3m��V@zsׅ����g@�*?��d�0�ce�:��=ҩs]X̸�;�t��G�BK��g���C��H7��{�Q��O32z�[,y�$�����Og��b������;�} iUi�ྮY܂"�2�̲��;%c�n��%�N҂1����{D��/����p�'@��{{�cDy�`Y&��e�>�1%{G����3�w�o�;�5�W�TC(��59|�E�N�q���o|�:��/�3�`#���`3�.���M[ċ����	�v�1�߽�����4����B�z<���Ի���C;+�[}ݤ���u�o:-�g�'�l���������w�GCu�kK
w}M�HI�j�e��G�H=��I����� T7ɑ4�6m�w��m�{hY�"q�r̫��7�����uH]M�{���{Y,���%���oJ��;74M���3F��9�y�3Q��uk��a��
�@� K:�]�z�n�s�e���a���CQ�kw�q���_�إ�y���B9�On�.?m�V2���ܫ�tP�e���0q��/����f�mR����Z^:�rz�&�H	}&��RoO���\f�Ȃ��_�{�>�?�ٙ�\Q�D����-K+�!��5-[}Z�V>Q��K��k�6�B����U�c:�c"�)�Z´��}+?���o�	��Z�7Ҵ¡�6��|%����������&�Cp�r)�:�;��t����Ÿ9��>DC��n�� {�Uz3�`Z��.�΢v�Ƴ���6ߟ��D�o\��r&������zdњ�D�UF�,c��ͪ��r��5`�U.0i(Y(��M����bϔ ��2�('l6�pM�e	1��Y�B�e�!��e
�Q�Xi[q1�l�A,�UD�V�ưf3�dY_`"��q,A��m�37�X]	](_[(��qn-���B�:(D���+3ի��RIr;���ۇ��?,�%�ſg�fZ:<���.�~)��^����1=7�� &�sia���O���Yw��!NVK��JI+�J�����inF���l���l�vD/�#�����C8ʟ��4�
(d"������J
Y}����iV�(8kj�>�E�&�w������mw84����p�;̂�;3+Ӡ��5E�s�T�2�@�������;~�7A�
SI��;�{=9��%���:-��r{�n���浭��N�e-�~.�H�m*��6�#��5Ѭ.
R9���R�©��+(&m�Ty2j�-|��8����Ս�Y�>Xb�}���K���
xUBx��[�յm_�( �y.Y3$�`o�P��)�����}C�ҡ�);�Ĵ ��WYK@^�KF���)x���=�k�Ln��͠%��8_>V��1��t��*�t���J�ڵiy5�駜�$b�18x���4�5�|�|����W�eK�
��770��r��t��j�U�9K�w]G�i,�@�kU�}�L�qJ�����TluV�8p��������g��ِ���S��jt�MG�|��g�4n�X�l���p��P��Ua�l|r�q<Ii�����4��W�E������q,��I&�6��Ǉ��h�O���W^�X���ܽ1P�h
#�D�/1y���;�>)c�o7�tޒAN�1��)�n�E�l0|�4Q��KPT�":�]x�x�zv�{���.r6����I��sGJp�)JOK����8J|�U~{�
]�m�3��qN���W'QR k����ڤ�����/L���cD�LeJ�BI!�p�}GH��C�h�#4����6�}yE'��m���ɐ,>��)x�*FA�������J�t�f:Bhx6� s�K[����dd!�c�l���T�T�S���6�J嫘�xO����1ʺ�k�vּ��f���C�g�s9i5x&��_v� �������8�]Y7K�9�uR���	���}�X鱧dj^����Ԉd@�!����b�5%���.nA���l�/��E�؎�-ȑT�#CFI	�5}ۥ�g��Z\Čhz�bE���J�́h�}��A��t���K�w�$D�\G�@�[p+�Q�4��Ĭx�`����o�ygT{.�4�ĝ� h�@�jӿP�,	5���/ښJ�V�1��g� ������g�B j8���X���to3��\�!+}�!ԭ��un�Sù�Qʹ��`�.�6i�\ŗsnO���|�;PjY���d�w�^��Br.�dr�y6�p�3�$�%��LiN��ӂ)�X��'$���|��w5�=UD�tT�c���sb�8˟3)�*=��Y�kH�T���n`��y�k^�/$]1=��{��)%�Z�7���4�x&��l�{���U��j\$	�����q�+E�輺�Nw�yL�/��2�z�J|r�=��!p(&����cG%��q���8�%�G��g��	,eO2��M�W`����H>l���tEզS��M��T&;�쇬S�?b���D���<�zcx��0D8�J���
��ğ����<U��c��s�F��L����p�A���X��{J�I��D=ٽn̈́�
b5W��Ǟ^�R���A)���A��})��k�L�(ҥ��������c��QA|�l��gq��Nq;�=��E���*k"
�6= @F}b��)z��}8��6�c���0��9;ٗ"�aN�!�ކ�DB�`')p��F�T�����pj�NaԤ�U�㐪�}�u�<kNX�Հ{����bHr�G��Z�PU� J2�O�d�h���������s�/�O�lݖ�@cb^M��ժ[�3�)e)><�b��W-�ϋ�Dנ�6&T��%Т����c1��B�w�T��x�_����ֲy�)�؏�~�/��TeW#f6���k�*�.S
G�0d����U��>;k���t��ʽe��;��Ϣ�橽�n�����%�M1y�'�>�iWqZP���%�H{o��mس�|Mr`���~��V�Uv�W�{OvhP�m!���Y3{(�@�G���Gn�.�?Ĳ�[ݜ><c#Q�Jf���g�_���d��5��pR!h���cf�D����#�E`Fl�m�X	5�����w9r*=5jQ�? ��V���)5 j���H����QW�����e��v]ݧ>9��&�}�De��|y�G�+r��)��#�_�.w���%�Vw���:���V�M�yhm)�̦��=�(�>�=�~����_�9Z0*#�Klַm���2n�o�m����Ԣ"���O�`m�9�(^���y��&<wJ螫�i.L="��Wk2_v#WJ*b��)o�L
t&g���db�a(C�3�îHN�r�1�F��e�9fEGr�ư���doʑ|�Ȑ�Xמ ,�j���jƺ�+IᎾa=���6N >u��/=t�{�[
/���4P�ܛ�Q��*,?=6���Xd
b3�7#�̲=�g[�����������ښ���>75�{)o�%T&h�0���^�$IY�M��_���:�����
��Y_0C|ث�e�/��7\�0Նt ��` ���3��l��!�ߴ1��%ы���~'w�g���C�{ ��w+`uK/S�^��T�,/!��y���ak�#���-E�19��<���k�����W�"ߦ��jMМ8pY�0��&��NO	�6!ܺf���j�C�y7Q��6� L��ƍ��AȠ��09]�auqIy`����U���ApK���^P��m���ǃ��c�����E�F����;�]�޽��t^��%�G^���,u�
����1@�gn�b�;%"A�����yvJ��gg�nG���t����y�Џ�R�����{K�)W�H�|=T�����S��6�КF� ��� ��[�wD1U��� 6Ll4k�Q��r��fL��qKK�+n5��i��[�	�|�Iu��vuM����Ea4��,�[!�p��+� �"�Q��:q�*6�uk��{�D�	�]V�q�����6#�����;��
XE�4r���dN�AO��G���*�<}(���wF��!Uw$�)�hs&ʩSQW�a����{h��ΐ/'��4��x�ը�T��|)UB{\�rE<M76��/�п%��⁘��/QI.��T�����1���W4�*Y�;"�@Z�����o��CZ�aI����E��v疝{r�����xr���{7ޤ�Y�tlL�G*Zg���Y��i^[ ���ǉ_�A%��x9���ϡ�r�
��Y��^��0�Y�ȘK@�_�p��Q]JG�b ��L�w{���K��zY-ҟ���F�7�\pޮs&�w&�� ��?���R�K|l&�I�v(����/�w��
ʳKƬ'�G�e�?��kv׆��������Ժ�O�v��ý�"�2�x��T��]�ۚ� ����ʞ8����n�`�n�B��T�t�vp�(sB��8�V�����ʞ�<u��H��/��璁���[Q�~ʳ"8��Q9�N:5[�l����M��ɛ�sݕ69������(�P\��M$"�������>�iU��H+�j�:�`�����6#\����Q����ʙ-̙!~p6�Ru���<�d=����k��=\��s �lFǵ��u��,͎쏠 �V�v���5�Wӆ�k=���8��{��=�I.h����@�!k)��yɷ@'te��V��D��B]��DR��Ήv�B��?���Z&�a�$�CXA�׋�D"�RH�Os�K�b�����ut��:�a.^ e vQ��m�����8���*�i��V�.Cr|!����bEWO�5�A��]p��s
5X̕���{W���Ja�Ĥ��9ߖ ���t�%�*�Rh6�*�'^�ij6�MS����0�g��&P��H�p2�@s�Y�P�w��A����?el��<���y��Z�.��N[k��B�naI(�H�J��Ū���^6 � S�ԘV�����`g���^+���_)��Q��Kx�O3|��N�~�9����>;Qѝ��/�Ual���}��Y�����=���}���$��k���+-]�zF�I�idz;�t���F8.���wX�rk����K���X[%g_[�M]h;�t��Ir��E��2HG៟��>��`0����A��c�����l-���DiHm�k���z�ey����J��D��8����3�K#�j����|���_�J{%�
,AU��%��ڀ��=�ą���AKQe����I�s�v~B��h���#��/ύ�G|:~��Y�ݠ���3�(r��6 �)��~P���y[nE�DP'i����P���<Z59 N\�O��W9l��~��"p���︜",=�Z��J�~�+0w��͕ZJ]ԭqDŵRJ�`��O���ih���Ә'�0(ml^3��EFѴ>��4�M���X��(����J��&���>�϶箳�%8��0�s7�|W���kR�c�Sp(�s��s��q�u�)�x�i�	Wv��]��!���`'��y:#�F��W�m\�K�u��tl��D��ͷU4�2L�;>