��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n����x>��r�_��S��7s�6J�t���/9���0Q�W����=b}T�-�uZ��)B=%�&�8|hnv��F�3�����V�}�ѧ4�B@F�jP �\��P�ο�����]��,p��2n�q?&���mGx�{#��@�9�_���nʠ� ��p��pJ�kA�9ӻJsk4���,�
9�y��w�e,��cS;����4P'7:O���w?�Y�o�������LǼ�l��Z%J�]�/�u7�(l	���l�\�Cod;��'<>w��1Ǳ|��e�0;�Nb����ʕ���Jm�'e�Ɂ�=��;���џ�!+=jR#�͔>9��u����V�ŨfA�.����D�[U��&;����L���w �L6�̤H ���DOc	��{X���-:J�v�<�(����ӳ�+ܢ��oFHMJ��Ww�ɖn03��V�|��{����A�c(G,�g%ʾ��Uf�@�$���Ŷ24�{4Q|*6�Y�0��AH7��<_rH(C��u`Cx�����<Q�����*���l���j��?�|��b���+m�/9\m �+9i	W�V�ڥA2��*.7����}������ն6�� �1z�N�\�<H�z�k3��9֯w�r*��ި�wa�W���t�|r�b�W��!cȐ݋&V+�R��l����*&N� �j�V,�.<=ncb�+[�/�$A�` ��~Y?��W��LB��B��]IGd@d�͐K���MV��� P��(�U(j���/֖.F�-Q:"�CC���ĺNݝ�_�<�y���c'U$��m�M�q�jlF�LX&Zۚ��}L��v{��S�n�3��`���ɭe:��^@��0���y�#����|�E9�̲�:?�`��n�D�՜7|7=d'�~�e��@�.�" -(W���H��d)_��wR�1�eP�ޫ�:jL���mh�
[gb�� @�;�d�)���΄�8�>�C�v�t~ݵ �K��5?j���쫚�IJY�_n��~9�a�ƙ�w�';J�.��{vQ�����~h�^�Q 1't�"�#>�I�d��� �{��({��A����S�n�y(��� ���B�^�i�ԒR3ؿ�~Yx�3�z��4�oz�x�ni�؇W�D�	���.�J�����#M�W��/8%V�-��d⮷1����2�9 ��.�E��7L=!j�˻\~�����rr�dڕ#,^d�/����z٫1i���܃���d�XJ��܍y�t��q�M�,e�7�ּ,�34��_�r�%�U�)�	&W)�	"�Q�HpS�_{#%�lD���DX�2!i�kiF��q�	�uY3�o�4
	z�<9>�@�U,��؋+�]�����4������*�/J_��췌whk3|S@��*��Z��,N����5���oaƽ+*�J�7��/�r���^�~���&�T��������a��̠�,�)c��ߧ|6�'�Ln�	s� 	z�1Ԣ��j�Ηo���M$��ǥ��B{d��w��e���&�ϐ%K����LF�4��`���2
1_�ݤ�{�L��˦]��6�6�����jNUM�i�L��HW-�i��8�u�b��.&�R�17Ա؞9KKmn�a8����C�zH�|;s#x�~�x�U�8��9V��Z��O��!탋����D��<f��gSA8ԆRso�^�'Ct�E^�NK�,�25�u��:��jNU�G� X�,��<$:=,I�ֶ�Ni1(:pNq�½�'�Y1os�G�3~c?4q�m4>���h;h6eY7�A�[f�V~K����F_s�\}�ꅢP�!�*�C��t�sv���� �5;~�1��\Ҫ¾��2EI�ֹ�v�Оe�Y��B����e���˓��;�k�Q1ګ�����Kklҵ��^�}X���)j൏=�z ������W�d�-��	����ߪ����eI�	7�4���n�GK��W���-rn�@X���-G��5(.˥��Vg���r��곇 k��ϲ%���6f�	Qӄ�G��|�24�.L�f�CW��파�	\�Иk���T�M�"R�W��MEP����}X<u 2���_�1���V��hK7&�A�s�p�VGv*;�a۔�0�<&ԙ6h�8���5p`�'�tN�t�xeA���vV��r�w
�
2~$�o��T�-����eV+U���P���+�{��A�cEi$+�5ixT�a���D06^,q� p��3f�|/)&!��Ĥn�{Y�6�*bm(Yr��������|�6��F&r���Y��#�p��(� �G����1�7l�ת�7��<����a~���|f� _YWq1�]��4�j��Gr�n��6����(���M�Ј�F��:�͛���ϱ�曍�0Q����
��Ot�T���,�NX7q���?����5�h�w<����[� �TcF`��$���@�izͦ��b>�뭥RΊ�Q��u}�����G�W���b2�_�@��F�l-?У���鷽�x��2�Bd�n����2�.�}S�^�h�^t�kӥ�8P]S/�d�MA�y�lI'���@I�)�-���[��8�)����B��~AL����L��xc,����Ҽ�ɪ����\��H_�|���ls"���.p�;T�6��RD[�����cx)���?��W+I�_Q�����lx[ �*��Z�[��o�D?�z���""?��g;[��=�Q~ha]�J�T��e7������ȡ� ��VP��b82��� >�^)����.��4�!2�l�X3W]�ڌ�oz�KA�--����2FiX�<|ey����uw�Z��a^�Q;/�"�����Hec|gJ�o?���� �<Yv�GV�#��uto��1k2j��Lﯼ}]�n�Y���SVL�Q����B�Q媺F7�6/��]�x�?�0�A#��rԩ�� w�Ig8@&�N���J�J��3��;H�f��(�������a�s���L�PO�S?���Q�r>�6Ց�8�U7t���Ӵ�.�]�ށg��&	0=-����\2:�>���A��eu�YU���=ϰ�L�]Z�(������c�X�XQ�f�M�ٻ�=���Czt�y�� ���L�_�;'��6$Ͽ��" ��	P֠9����.o��oŀCP���+�cɖ@�s�r_���Щ�`>8ͻ��ϗnW��N�U&��CxqQ��_��P�D%�nG�(,vG�����H)��	?�d6�C\k�s9�n��j�*!�r�|�m��8��N0���%�J֤�(��E�/z���Ҹ�jK�q�U73G��Jc����0DP�N$J@���WRn~�2��"#~�{c���Wx������Q|#��e�8���[�8��������5����^���q:a�/�4���E�sl�N�Uf�ۧ��t�T���ck��ph�0ɺVxj���^��M�Rn�Ű���W;�����S�e����ؐ��S�a�7��g�����c�l��r�`M���~��,��J,5��L������G�G��Q*)���.d��{L$U�^�ܻ8���ˑ?��y'����Ӧ���U����-g}�O'��t��8��0}�1��^t\��W+'q�^zn��ea�����-tO��]cu�����B�����ܠo1����	���[��Kq�x7��r�z��̧ޣ �ʘɑ97��w�+�so28Wt+�D�Q�A+K�fó)��v(T��p7׈��wS*��Swvڸ|dB�W�]i���!c�΅Mj<�<�;�[��Mf�M8.�+tW:	������B���:��f�g_&������ v٫��멨�AA�� Y���ޥ�'E�cBc��5A|	0+�;J��Q���9�����&��s���� R/�%�{�v�L�;��{�W��t�_���g�����n���I6�W�Z4������Կ�`Qs��B���FD���s����mB��QOZW3�b���cP�+P@-�D�@G������=�S/]^�}Б���$����-?�X���:�Ci>zL���t�
���4��ߧ<y���)��~5����-;_�4�A�A�-NA�m���ތ*%���*+)>.��i��@	NNo��s��9,N�K�㐠�ڻ<�,�I��T�{V ]�'#R� y���s�K�u^Z8M�{̝ļ�0^ITy��%�}���{"�*!�G��\��[���@B�U�M+tk���O���R�0���|a��Yn@n��U����T��h xBPQ2yG̫v�uc"W�0��`P񰋱5����D;H*k�)�+FUڑS����Aƒ���X?�T��ʁ,L"�ݏvlk�e5�O5�B�����bpB�S��M�I�Z2��&�I�hf\eŢ���J�Hws�^d��G��xk�w�� 3i��,�B�7Z�P'8�67�av�O=��I+�W�8XM�3�_7�Ys�^��Ǆк*Ӹ�S`�mA�Uz�)��8�y*���<t�6/�|�QH'C⶛�(e��ƭ̇s?�
�$2��W�$��dY��/w��cr����@*��q�?���r8=R%�s�bF�~?�-c���y�L̗ەͭ���(�F��� =��U��/W�B�W��&�)�@���y����:Q��������v��Q"�Z��r'?*Q��Ȅ��Ll���n���D�dΠ�"� 6aI��)��� h�*���[L,
��L��4�W�`���I*���a�8�s�Ws0�@�=�K/W��ኸ���_�Hնd�I�aD��iߦ��
j��9��+6jy���x������5<�������E��x��M:���N�/~����\��\[w�:�ٙA/�����z�,�zvp&]���U�j�����>���S'��U�����h�'���= ~o�E�,|��}���
��|��ڜ.��В��H\�����ͫHs��`ug��C_��O�09�>D~�!N�X�SoC��*�թ�oR�fо��f߽J<�[K�W@>�����E���j��X�dલ5��pBݦ�w���㥟.þ�X��5¹�K�4�}�e�MH�Üu��\EI��U���8@�=VX�����s�ާ�G��\�`�W�U��+4b��wp�N9YD�����qNY�6���� �Onʶ*=���p�M�|��
����/�� ��H����Y�����m��R�W�/�h�Es��7��n�����we�3v<��:�<R�!�S�y#
WJb\9�2%}s��瑬�}/�>����T�H ҫ�ٟ�(l�c�q��(k���7����y������y��Ej;�2@�/�y��t��%!��^m9�ŉ]��C�܇���1q���_����������N����d��+��n3p!�ڡ@��ȡ������+kn�-[��kz��:I��$�xd��)�h���IӃ�P��d�:����%�%��O2<��1����0EW�]��=�S{;p�+	��@�\H�i\P-Yk��8!E[�r���!Na
�0��l6~t�tx���@�bٙIqX�@��}y��G��O��mޛ�#	%��h4�m�A^��LE·%<��y�z��+�t��b���T!�㶟�����!���܆K��<J��}	#hhwX�����;��9�0c�9�F�{7�m������н��,�JBUX��P��w��P�p
������*1L_��gu} ����K1ɯm���k���\�f�P 9��{��h����)	��yx�~`�2�;n��өb7�X���&G��L��G����aT��d.X�dA�̯�I&�����D�4o25'0��ޮa�bn�pڡ�]�,������C�!3��o���c�o���������%��ߜ�#ugxŦfMh�T��[�0�?�ܨ��Q��E�5�����$���3��A|�jȊ�d�\<2Dd߉�Zt30�䬺�X�$/^������;����
`j���"���©���ȬY�L�$���;ꚉ����^���>�|t�i
\�J� U���Ρ�K��&u,d���� G)E�CL��HO7�{<��K���!��H��z��	���Z��ј�_�-�.�ɷ\�mu\
:�ͅ�J<�,�ٛ�7;��t`8�X������`��g��ff��`��Q���8A|�y9�W����틼~���p{_���os_	p/�[��l7��ښ���"4U�^�������gۛPD�U2"ur�!��=͚"�K7�����t^�b�rƷ�aHM��t�Xu��������������D��ڝN��؂�\��+��<��q}�^̎���oa��D���j#����dSr��^�EȻ=�cy^��[�;M&�+3h����m�Lڰ.��{�C'�9�	Y���J�C��R�{d��p�K�)[5�
�t4��^�τ3{����8p�;�$㧌��v�l��� �4����,��B�\݁4%Zd�p����TcI�K�L�a�߶��jsڌ�]D1C����x��y
=	GLq�믤ws�=�:�0`�E��}����^����=�oK���d�Ef����O@���л��R�aׯ��� ��fyEԽ��F@��ku?5co+1�E/�U�N����z+x�1#�!z��6�����t�u����\t@0LL�Ȫ#C�O��L'���&B�K$��5�A�*�����=�++��&�������)�/�����J};��x���[����O@j0B��"����)6<�s�j��j�{�3e��}����'��|�q��&#6�_��G��}4'�W;C��4�"�뚟Ĉ�L��3i�.MQ��hr=�����pLC�4��A��e�vG���Fȏa%. =7C���L0jySNݡ)�&�iZ�^,e���:7�է�b�����+V֦��l+�M2d���J#O+:'�M{��O�|*��'0�A�[��r�S3!h�"s���K\T_{b 0�j_����7n��
B�(=�yS�uH��#�_	{ث�wu��}����9?���у��5���
┳�A�sұ-(�/���@[���x�IO�+�3K�2���;w4�P`w;� �q	�"�'��G��~e!a{� �#��͞��y���b�g`)�B��AlF�㦉_�zҜ�_[Y��D�*��R^���9�lBR"�ŏ��ҕ.�P}}�]8����DE�C��J�O
i�CSc\�e��]U�5����U�����|(U�Cߝo�<'\��G�����OН�Y����7�"���״�p�qi�X��ƒf'�J��X{��s�	΋���c�W?�T�����e��gX	�C��@o�!u�j*�^-�կb�p�I���䛻]�����@J+N��{sR鑽��F� � �h��K�^p���<4fȥm�[�G��	���<��h��k���qf��q����+��?~U��э�ד2���c��=	&���F�Κ`Z�NP3�9�m���{�/��[p(o�Zu���C�V!�h�Q�n��x�?���|+�T8[&cםa�[{@�'G�.�M���}��ؐ�fH��Ɔ��_��Y�U�C��Ϋ�#���ΜY� �z~��]�cm��X�ׁ��ѷY��<��*!�OTP ����.�F�~0�6B�cm.ý���K����g;��/�RP�������p{0��[��I�,��GH�~�V���2)�g�5��hAU��R�È�قC
`��P!:i��`�^��L-�<��Z��B������ߙ���[⽓<s%��5�_ߌ{� x�,R�*fVD��>�%k��@��"*.6���T!����~Lg�?1�Upu����Qs)�{�\��v�>U�c�2��BV��~�|���Y����t`��:g��}W���U��Z�M�ڙL��o�n�_�+@�p$�3�~��s>E��[.Y2Dd�y
����p�6���c�`�2Qb�^�<��P����l�Hx�C�E��OPN�d�u�(���:�g�����L����+��:�rZܜ���8,݊�ے�X����1Q-%!Brz��6��I��a=��Z= �X��r$� �&Gѫ:��k�(��C?�ӌ�ta�G�
�M)�y���0C(պㅖ�`Wа�aRg/��b@HU�ѡN-��٦.�����a��W'�V<נ�"1���,m��7��>��t�Q��H�.Fԟ�_���g)�b>Wݪ�_)6�ok}y�
�u7ѩZ/]�%�|s�ɍ�/r_�=n~ ��'�M�֎�p���y�T�����e�,�h��_��ξ�v�rt�#1P<v(3����Kiݗr�f�]F9�&x��j����S�}81ʃdEN�����aUWn��>7l�K�{@L,,�#�ݟ��>%�����r-e̜���V�nS�M���P����{���e c�G{xNA�����t����Jɕ��e�q{�����?�|�L#8��7p�Lâ�I-W���<�._[�.�,y�'I�T�>S�~�V�#�n���rV���&��i��0�9�"�e>ָ.9p�	��p>�� �r[ڮ�%�/1�M��y�0��Q��Љ^p'���m��������lG�)��5�sE$!}cΰT��n��:CP�=4�o��iI�����L���?��a�X�KI�rc���wt
c��a0(-���^Y���*,�;��sl��c��O�ዳ����5�	�	'��9��^�|K?�ǽ������VB�$�T�Suv*,�����=�'��-����Q�~L��Bt��#,��O�3�)�_���!휩��TO�!�s�����FS��<P�m�ǖ��Cx�~�|Hk���Nf�m��cO��@o?.%� T
&6k���|,�\�����H�~{��>�[��>�!��"���:dS*�����K�C4�&��F��-%YQ|t f��c�Р�`[U�j�̈́,R�h�w۹�2Z��⴯�wt.ջ��P�I��6�#DI��P%��=vkKo6vrp�"�^�^�R�`]v��Ԋ���U�Og�)�Mqn��%�Bg�;;<��_���q��}`,�µ'X���>e�����#��a��X��8b�5a��~]�2
�)7�����,fd�C�>�e(Y�b[�帑�BA`Dt��VQ��b��������hi�S;&�p�X�c�C������my�~��)�����n9��:��l�ڿ�;�(K�ѝ[�% ��7���D�i�Ek �Nȴ�U�oL����c���z�>��" ٺ|�U6�K��H8��,�h�;O��W|�Ńp�y?�qo����toa�\��[�������NjO��n9 Q��\Y<�y,��!�Ą*���g�f��N�j^�Cp�-��g�wN��d�$�G;w�$�p�+�q��K���*y�X��AxGp���m��0����Ў�|��9�#��-�����XH�>�	�\�-�SMH�p���`T�gN�5y���u��_��G����w���;6�MV�C&q�u�nY_؞p	�L�O��K�h�� V�	ϫu�NS�&J?�Z�� ��Hk|\9�~��=�@�J��_Z�H�U'�o���"�� f�&�j1@p�<r>�-H���	�Tl���D�A���US�1���W�R�{������ٕ�Ԅ���"!��Pkȹ��\Pp���J��j&z|��^x<+"]�@`9u@�<�A�~4T��Ҡi�ܣ7)�pk��롶U�NCCHNebOO}�5������_۽�Hy����M 5���_�%�
��!�Zܑjn�ؑ�~ ��	���>�=��H��e�˨heI&~���+�Q�����.Ҿ������{��-��@N�ѶT��)z>�>k�AJ�(5��V��st���]UU��(�pJ�5�kB����|;3b()�~S/oE}h�·/�;pȤ(��P�����ԫ�������6A�!c�4v:�J���
�;��9Nk#���Xf����� ejd"�b*�3kZ蠻�Utl�^Ӽ�>��u"�����!ˇR;�>֎[���H ����x�`�!��s>�wЪ������k�h%^+ZW�����a�u,|f�q'L�}�btR�=��Z)N�]1`P7�|�v�!���@�&k�gH�"� �
r0&Ta����FQ��O0�.8����WQs�hR���+H^�{@�},�";J �����ܚ�0�����V���< %��Mx]k�1��7��	��DߓQZP>b�B����t��4�\B7'�>-b��h�8,��	� ���,̫\�nER��G%AY��]lэ+J��f�#���=r،t���y3w�3/�FW��+:F�
ա�G��@�w��)l�9������ ���A��m��(�QK>'���.�4���+t~*ȷn�n���˗1���b���
B���IA�myn��i��22�ȩ��e�+R_��(��?�}�ʖz�UwX�������e����0�7����-�goe�3TZP�**��дX��E�&���e� ���S	K�(s
9��!�%|-X��i���hH��"����ࢁ�Ya4\t����j4�D��W*�3j~|�e��b����4�18n?����p nf����j�2X�H����<�����'[��SC3���3���hF���~���@�H�\�sy�A��v^w� Q����	�#��'巽?�B�|��(�q��Rvl���+r��ߊ����(���r_�Y۾� p ��(�=`����W��S-#��quq�fN��(8�M�+q!] sOr��I��ޫ9�8����5w�\�a��L��-����/Ҥ��k0M�H�����ȕ����=5��Xm���s�A&[}['ٮ'9���^�q[PXA�ϺHR���~���G�
˂>�5b���f�)�R��>1�x�{�;�ߵ�I��Ur.�����E�.Ї�����L�"���`�@���Rh�]ǁ���E��1�@f˷ߤ�����`��y�����G�Ϙ�?T4
�<�kװ��O$����qr�Z��:�H�~��ꔈd���bc����!���/��&Qb>��S��9(�N�ߧU
�"�ր� ��1��@��iH-p�[��(?�m\��>��*�4ns[e��hWK�E�2�E'��K��m�7����!��O<� �iA�P,�����_��,�fu �����3Rl�r헗�X���Ɔ�L+�o ����;�$|!�����I���C��t��mC�������㯩���w���8~�����a!dj&
���o��V��Me�IcM�W�����;Ss��S� �<E���#��0
���鹯�j���k�2�2Hn��΂ǯnB�9����դ^C&+�:�?��侸�h{�+5���t_\�w�S��2)���؈f���Q��v�IGj;O��hOz��U���&xM� ̦@�c^jCh1�ͽ���޾��%�@'�b�J-uR�����w�,�0R�$� ��:>��D����w��7]j��9��C�D�%�E��K%���~�~Ma!|��]�@�Hto�\�����&�O�Zme��~���FP�"Y��C�~4R���D>f'�8~�~��e�i�2�3PI�u�&�1Y��1����od[nL�Rq�*΍��щ.CO�����bh��x��EUI֑sG�5/��qX��Aa}L��P'���,_�|N2��=йn_b=O�rn<�݇5��Iq�e�0z=�=��ۘUW�}b��`���.P�0�M���KP�!��iO�����VB͙�V��_kY��A�d�k�R� ����Ikh!�tOuc��P�j#Y�GWc����g��q��E����f|�ZWM�6�����z֢��h���E��ϩ-tt��ȇ����lΒ�l��8�I�r�r�v��#WJhmM<�?OSS�B�w�	���p���&�WIPEqM����i���h1���IVMO�,���%U]��U��h�Krb��
�r�L�z����gE8�������˙��Nev!'e�$e���nF�7O#��h����Hi�4�%�v��?ff��������oxH5�Fm���݃�hX�H57�t�h��q$ ,E�9c}H�N��r՗t�+P&^���bWV�~{Y	�՜��#�Q:l_�jx��0�ȫ���{�.(��,� ��N�����~�D�;�l0�Z�ގ�8���C���$=x���¶��L�?U���|���J�8����A�b�4��ta<L�W(�A��>XQL۟R��(7ߡ�L��0�+����O�À��$'�]�"FH���Ϧ��eh�L�^���>�9�T�5�s����ӹ��&�>�(�LGL&#BD��"4)۴�5g��Dz����MgO�����t��^OŌK� 9d��ɥ�\5��F�Ka���+>1��t���*�t�k ���o_pOEr�%���Fh�AF�����%�|��'�`+%�Z��R�P`���&��1�8��
�Ѱ��G����?cTto4.Pd�o���[w��� +���ܫ�?-:7т�^E���I�cC>��@�Rk����?k]��(���ul'��? �Wc�q�p�}-d���q#$,by�f5\A��>�@�$��-�ğ��(��A�/ޑk�oÞo4�'!LA^��Mf�َ�w�����C~��ʱ��YS `�b] �Pb�R��#^���JB��fqm�&Os7yk��/�~�z�Z�����$����]E�'�qw,H���hi�`/�=���L�qD#�~�;@�B�{7i�R=^��ص��ȳq&�+Szo��7-*��N:���[��zjK��h �׶�����9����|^���:��]D������_x���Lx�1q*l���Y7���bg������Wu+�z�Jd6�"��c��į`K.B��2�b�0Ȩ[�b�t�����5�Esoh��blFl��ȩ�z��H�:%"��� �-��R܃fj	����jb���4!;��ס�RN|�e���:/}�dؐs-�s��OUu�·�Lw$�����q��~��"�i����
v&� -�1Ί V�{^�M	�s'�T��+�	6�h��s`��?SP�����)+�Nս=�y���M�Js�gL�}C�	b�/�	aW�6��6�h�ŗI�±��:Z[���T���DU)���z�>��w6����@���j���;]��=9
=ڝD,�Y�'j:�������KS4F�e�-���?�J�t��8�%h�'[���
�V!���0 ���S�N��M���u��bꚤ����ݕ���J�(!��k6w���\/�he��o�b0!�}T�g�(��~Jee��05gQ��i!��_!W^&-�i��\
�o8��%<�D�g{�#O��9P���\�n��	g����ߥ|�����a������[��M���[������v��8@�U_�9���&�}9اm�j�}8�Pu�T�n:`}����-�j��4ꃺ�c �S$�\�ĺB�[{��yP��ʦ5p>w�Y��	�]m�>����Ҕ^(U%�y/��E���	S���LY]�	m�T��ލE�e*jc\Q�bP������.t�v�-Z��i���/��yV`�o�Y�<F�X��!�͵�dc�VN-M+/��bm����Tw%R��a��Wp01����nuKq��O-���[�$~���c�'e�w���,�ì4�"<�(<���z �؂�4��g�&#��p��]T��r�g]B�Y�3���9���(�n���x�$H����-W:��~����/��v��r�<�\��]����*�jj���Z��ZD�'�pWƇ���o��/�gL�7X�����	SJ��m�.br���$F��o��g±-B309e�=W�v�LFt@Yf�?|ͱ�s���C�B 'v�[7.#K+0]�vZ��P�l�d����]���
E"~��} �[Q�g[��q��QN�},������!�KL(Z�n�a4�p��s>O��;��t��v������0���9L�ŭ��e���M}�p�a�*�|��8�O�j��fߜ,�V��$�������L��N����K9lq��Eԉ�	A��?����g1���Yi�"'*�*E�;/W��v�O*`����	f��(]�Zͻ��}��?���4� c�YA�q�]�"kˑT�6Z�:�?�6�W��~�i�l��
�O0��D�@�D;�ܝ�F�hB��L�j)�T��$�@�w�VH���3�i��t2����Q�ÏxK���_k��+k��0�lW����wܽ�Ш�d��/��d�� �(���L���OےK3�]k]ge��r��1�&S�+$����Ɣ)J�M�]�DB����n� �t�h�5��Ir:�]<Ԅ��L�GORR�:ғ8�M~��Q��)q�w���	����ѕ[!�+H�DRw�',f���� 7�;;�o�/ZJD�֎��uؐ��69[�(`&8�� ��^2m6��m�T�po��2��oq��}�W��lF;vXXE��o-f��?��O���|C���}oH�-���N�^�X&p�א�Oz���eX;�8AQg�Zj��-��۝.��M�T��v�r+I��-\ˀm�D��T���s�Q��
.��0�� W߉�F�X;�����X�M�_<��sp��U�eḿ�b{Z�&9�YSw�W��B`y���%��Z3?��bj=�*��	���m�~#+K�>�ߝ;j�Yޭ�*cK	/������r��[�7�
�a`+:Z�d5<��?��՚N#���y��vO�=���V�����Ɉ��g��zMg���K��Gu�!�LX�g*¦��q� ��A����Wt���ꃶO�Lzhۣg���stK�p6��P�d,`Ԛ�����Ѧy�����$�a���G1�1�V�@��^(��i�\ LX��������R(]vm�]�_��^���vm��z�9{�M,X~�����D����cA���j�Oo�-5o>�K=}���lsU�����C��Y}Au�H@楶����W�i\QZ=C���	��z�UJ)�*<���N�-kF�����I�2֮�.k�^}H���'� @�D��$ȒJ��|y���䷓Q�d/v�V����ևݩLs�����\蔁i3�Y�T�Վ��d��k�ck��2�S�&�]�t_��2�c,%����b��E�{�����Վ���Z���h��RX
��TtN�����s�r]f��E��Y!��X�mU���Ƭ&#��
0�;�u��ٍʞ�d�;E���RЪ��e� P�m�#4HOa%�[��w���P6�C��q��+.��>x�I��Ҕ6�@�Y�mq������-i���&��t�&�9��:������v�PQƍ-��N@]1����+����N�"�˰yoe����. ѐϪ��50!6Uv�p��e]Y|h-���x_���\g�J���s`.�ϐ��i��%��lG�6+A�P�4G-�g�فҒ�c�!;1��U#Du�MB�3@r���~ �=,��fr �:�-����붢xY熄��k�����1��w��y�Y܃(�ө�rvG�(IJ�9���^?�ѓ%���4�+6,�%�����Y��Jk�W"K�WCN@櫾�f�Bfi�Ѐ�P��<��;0��2љ�ç;8�n�!y��MQ�";)��{|zi0)��̱�.Z>r�d��`	�C�+�&�:t��p�m\�2uFzQ�����b�C� ���[�<����:�ϻ� �4����-�䂪xz���*�T8�\"1��<L����u ���$�7�Y��������?����U���w�e��d7/鐵��
����#ڸ�ǟ;OL��/�)Bu�qx��Bv��uc�C�ۛ�S���t:�+,a�3:g��)����gێ�c�BF�B�Du!�����nEgC���y���1̆'9��%h�݅��OGG��!�C��?F$����W
Iإ?ɕq������[���2��=��jE��\j��jc���\/8t ���O�x3�녨�u�}$�+�:l"��:k��f�29������0�q�1�$��\�X�*���`�����9>�`M�'���g���.�"�˨�6 e??
�Omkl��9��.����s@�m�y}2��X~Y���B�H��Օ[���)�vW'm�#�r�I@1;�ja���8�|�92�.ZH�q�7�ޭZn�^��"&��p
=�d� �J%ZRT9Z? ��L������8����Zo2$�Ѧ&^��TG�l3"#`ֈ����)5��摸��C9��5�7�)�M�@B ̋?H1�\������+hB֥�5"P}j�k�Р�.B�]R��Z\(ھ:c������Q�Ų;�\�'�$Q��-?�)���Oih�ar��,Ǌz;*�|�,Dꍚ.(��>Hd-���o�׿O�\���О�� ́U'{��OҦ/�P$:}�J"�ϒ���L��j��snr���%��&)�+�Z��O���j�n=+K�O�^��>�ז>ۮ�	�R�92�MUp��m����I�����{�pC�;�BZFZ��b�豁�s����$y��k��ې�	Q&�������,��z��8��[���j���84*0�M	��zX;F�a�&������`;�$���W��A�tVH�Mk�E�2�#_��Hԧ ��ͮQ���!�L(�:XZ��f3.]�;�!~�`E1�8���q
󘑗4�;�q5���G����/���fҊ��ksV_Q�k�s�D�-Ϸ��-������ 'G����4$�S��B�L��td�&U�� F5�jԘ.�d#qp��Q���#�W����:)'橖mvم	b�o��,��J&%�3�,
�,LRK�$ݚCb&��v�Dy�K��_#`�&2 ��\f��vF�4��Z��qХ۵7q�|,.VC�����e��pcn�ջYK��Ƈy��A̻/�W}�:QM	��ub�P�ų�qV�w=�]x{)0KQ2$�>.V�#I��#LA6�D��,��%�u���6g�gϱj�q%VH��ʋ4���wmޛ���]�`������z���|e�����ox�ʅα��e����'`�u�� F�9�G�+}ڵf����m�1<�X�g���N��ꏿ�b�0FLl���4J�G\4rPx��qX� V�H�.���]�b��Q�9�}���������(��p�t��QaTv'�R����xV]�����Md�y�3�.V��y���dQ�F?���J"A��JEΨ��f��z���XJ�8�u��8l*�QO��u�	?�:���˃K��BT��d�G���Ng��N�� 7LA�8+�ł @r��B���\�����1�k�$|�5l����$v�����^Mdrȡd�e��,m�7l��ʾ�-SR����B���|�\,��x)�'�kh�9�k�W��vYb@�P[�rW���|~w�<RS�UH7=�����)
�T� uO�����e�����s�8`�v3�Mx�+3�}i
h�� A����|W���;F�����	,'��i<Z�o�.�2�����9����1H��쯍#AV�%av�8t�`�]G��0"=�J���~����a>l�Bu����&�uX
��,J����c
�H�v팕�ll<Z���J�N�)~A�@�+O3&����,�h�T����D�]P�ܗ�oʩ>c\W��V�U��;;�����Z?S����Ϫvi�H+W�Gj�[Q�1��r�T�v���G�眯�Ÿ����c��\_�o�$1+����R�*��^`����P��fR�sN!d����^��~[7��s��z 9ZYQ��7kxc�?��ݍ:n��\
��*k�:�1��i����t�%~��*�j)��|�r��C?�a��{Q����#�D�VI�@�NZ|v�ќ��S�F�Q�C�8�����>����3���dc�_����n��ll(��������>Գb���1Tc�V�;��9��Z�����o3�T����~��,�v����G(�-Z:��9��5��7�8$)�e�<��f	�
�X)��z���E3#0���ռ�q�N���vf��X�VC�Ӑ�h�h(a��6�AF ��w1X�U�� G�;�� �哚�U���_|G�-�{#��k�>4�NE뙄,Bi�&c]~EP��^:*!u{�I�I����,ڻ��3�� �d�<T)W8kM��vO&� �+U�rA��Hj�E[�x���h�WX{��۹�Q�)<��(ܑ�!1���> ��H�V�%�Y�ab O�-RL�@�iu��g�l�����B*���jt٬��,�4����}�Jʫ7]l��ZR�aD���R����&��<~<I��ֵa숇Cp���� !L��nJ����"!��\�pUi�>�b��`7/]p;�̽��[��Q�����6�����%K�p� ���#T�4
x�8c����ȵ�)���rgЄ�~1g[*���V\�~�@��P�Yyq��*_ģm���R�8�S$��Z�"O8ч��I.�Q�W�q�ucS�D�H���y���I�#�MT�7���4#�	�u(g��~G��k�#�a�]IY����^tfs�I��B��
{�O��g�|����w�j�vJt���؃G[x� EF�n�*"���2�{�Mh���@�/?(C[j��!OU�y�}�E���F�'�߾���3�B�E���9�O?;F� 
֚�����**x��i�:N�Z�r[��w�V�=�ϰ	V��t~�ÀǶ
��S�� �੃��Mz|�ʃ<`�Q�?�ʡg+E�W_4'�|��g>Vdkuܴ��W�-B�bn:�(�c����?TBki7�U�*�`�a��E���R�N�6������]�ժX�Ҭe.mU��K1��1��q�0��%��<D��i��2�,\,O�r`���ЫN�m�?s�,���A�=e���;��2g�J�v��P/b���c��۲���G�@���$	@g�*��y��9�d��L��rm
er�E����\pM'6�d���}����� (�Ph�X��+^T��ƞ�;���R@�u��.�1�;��"�F��Y��	 w?���K�QWY+&�>H�2L�ܳYF��W!���`�N�lEm���D��%69��=Y����e����`~�cadѱ�Uټ@G-�{����P�ş�8K��x��e��
�,��V#�#�>�1�nD�=�H&�d-�����UVXAKxaS���/��^EZ��Q9�	�si5v
лӌ�Y�J��v`�ж-KW��o;�lb1[��t��
 ��*�e����)b�)�`��8�ڰ7ߨ���Rk�b��]R��TJDW��˷�L�����	u�Eo���i�,
lb�R7�gw4�&�,�B�v��E�D ��j����M��cR��6)�	枈kf�F&��8#�2�ϢfG��ғw�}�[�E�f�q�a,�>��+qL`����	iB�h'�)OԞ�O�-�4h#��H��b'sO~��E/�E��x���(��������iʝ<�l�	K�}����ub��T��AI�H���6
`b��Ƽ�u�#��0���g<��h�66S*=�l6�1|��ObB�����<����!}&�$L�ǴM>�@�;RO��߫J�~IW*�&9�n&�꧃Ae({�]��Z�nUO�-f*�Adt	zs����X���8�
���b�%䎀:�X��A�=[˦d�P[lb�����8����D�^N淋�3�W�S;��)������;X���2�.X�6	#�K_�ن71I/���-H�G����/U�ٛ�u�;�~���(��O�j*rЃ�Sd��:>���f��K����[xD�!Q֙[�k�K��D4Q�x"}�%��`O^ �M�fa�wõ�z�<�^���Kc�9 V&P����1q�îN�LV�u�]Q�o�A%B���l���F�Q>՘������*()mcV^�#�[�\X4��e���2��HZ��&�Ñ�NG�t\�Tgׅ&c�</��uҪI ��[�>���I��ke�Ε�ޝ& !���:���}Ԡ���R���������KT�/��A3�����kD�/������̪Í�����;v���j�wJV�s��O��$�m���1�#Jл~���\:�3�m0e�j�iZ�>����{Ci�9]�|I���D�%�k-u��)����u����BS�]B�|M7֣qUU�0�I^H�<eօM��m8�=/�|
���[Ο�G7��A��+JwZ��ma�D6b���:$�2��W �����b�H��D��8l��%onh����;n����]��S� 5��>U���Ĩ��`N�h�_}�h?�����'������廉�h����Ω�5����z��m�R�B�'cp
1�gN��Cn����kD���-.�@�ܕBS�hK�s`������*�б���i��s��7�Qt���f	#�X��k�G��[��8��Q5 �X�����Y��="���ج|��9���顭��F���'=>�-@0��zb��@���L��N	��z�	`X�F�?0s�xM�)��Ⱥ�*2K�Q���;$zv �oY�T�yY�σc@��-�)�3���%�h?�6���I����V? j������Č�^�D�@adD!�n-r��1(Zpo�����oW�ϰ��*�����������!U�)�0��$��z�C.~�~�r�ߝ
��saURT��Ѯ�_���g�PKF�n��Ym�G (��	�5	�Yn��V��ƷL�ѥU����x�}S_�]%s�>��/��@���9Z�x��5��>�J��l��+e��l�p�!|���&��x	�t�;﹐Je-]�ދ��w�W$���+c�9�>D���ϕk[�%o��F��`��m�ٽTʊa;�RSl���]4E�������G�,����U��A? ��
f��CM�n��:���p���l���C]J�����8�_5q��1>�@�
x��=����<�g�*���]�S+�zdO�M4<��$�(o��Nl���]�c�ӫ�r�Fd�c���'��g�,��g�x��[ufZ֯m���ӿ��J�c�V$��`s�1J�c�m������]Q�+�/��ۦ\$˂�S.=����5L�r�[�@��a_������eA �'����Bz4[�|c��:� y�7�M@�D;�-�
�!�"+�� cG��肎@��X�4�4�̱�<}��S��<1 ?۪.�?_�M
�
a@x4��X:��UE0Y������g����]I����kO�S�
�b!�X�XW��ca���5"NɎ��hP��8���g�>5o ���twkT2��:6�#��l?�Sɍ�D�S��ܴ�1/�Bj*��X%���X��N���F��p*JԂ)�h�&`���EXf�>�2t�\g����c��BԬ� ��yV6������x&��M{d�Ӡ~��g�y�����(W>��%g�#1±�8Tߙ9mu��B��JW���2���ŽT��@!�6�54�����2�
�7 �T�Oy�(Ի��:�3�	�2�_-��h���N���#~���QO�M�7�%~S�IO��I2��	�;��-�f�s�11���Q�8�R�b%� {e@��X�#�xW�����@z7�z��u��Ʃ��Z�s��i���+�}h�^�PmZz���:a����K �-�1Lb`[0+�ٱ6��H�47�	�DЍ}�(�~|�Z�|���V����)pO}̠������P'i�]��j�D�V�s��v5���ψA�(��|�̉�{,1���3����݆w��9��ُ�qX��J����J�n���O��̨��yVʱ5K(�A
���)�J�d�`�� ��#� z�؈>p�N�5U�
�U"�[�y�S�F��4�u��s(���J�(N\q�I� ��&U�����[���1ia֊<���$W �3������dN��|��z��҂E� ha��:t�f
#�$�L <�}M��$L�gq�݇���JV��n��/OCuZ����t6��E��Tn�:�]ű`U#4;���;`�D��>�1ɤ�҆�B�)!�K��^�=/��OH��L�����t�Vg�D�i��*�rf�D�>�:������̣t��R޺M�2���:�:�Ɓ<@Y��E�l�{X�5���4��e���,9.nv=(3a�Z��2h�Za)��&��)bZA��6�(Ky)p���=^�ς�ujٙ��m�6H�F�γm���JUh��.߆R	A��Hx:�"|�	j�&�eI�;I�����yr���[,x�i�+�V��7켶+�U��y�!��1 ������GHg;�ge��.K��OX�@I�ҜM�l��U3�X|��%�E���K��=3��k��E�d��$ |���g�}���ՉD���9��gJ(�	�b2 ��ԅRp��! 	<9.��Hz�R�+n��Cm��^����mu�#M����p�#����R��3k<<��=�\s:��]�,Z�<����ST�U�,
B	�\5p����w�z/��*�	Mjz]#g�Ϻ<��k���ˊ����Hpw����o����3�����7�u��^	B��1T8$���M=��}�E���w���S5�9]�%�:O	J�����|6P�ґ<*8��`ݖ
�'�Q	-�;���M�pŧ|[�&�ሞ���@u%����$�	=z	!b�N�M��J֕�23�d�\�F��t
��u�t�K�s5�ZN�;��	�g(�!q���y6���l(\9��(���g��:/�䫗�Q�gz�5f��6A/S�	�?6=5��$D�$�d�Oy��]�f<��/�5���p7�*W��tFˇ?<S[�N��#^�A��#C^��qo�W��
��`��|}�����S �ٟ��O�h���O����b��PT}B4HE]���8c���K��:��^GG�q���˧�j���G 4�i�pB��)�?{'����06)�$�UK2�Ë�i��u�����>�z���N�V�c>�����ܕ�Ɩ6r������M��n� �Bg�d�4B� S�����	
��E�uD��X۪�*��{�����(B-��`�-!{کv=��E���L�Ne�3D�Yl����&����ko�H<��;68՟��%������Nd:�����]�!4J���/�ۙ�D�������+B̉�|;R1pE��AI(�zp񷌊�C�Ntz@H���'H���ډ����:GfA��Ǩ��B:��zte���uo�p���1�KR}x�5���gݯ�]�0_z��������G���z�J}�c�#<�=v�h*�h��E
�}O�aN�C�s2�.����v�A���6� i��S��57p�j���ܳ^
Y&[�����eS=Y+ &�?"3��4����s"!�S�έ�wz8����5�����Z��Ce��z�pwv�8j/���i���*���Å_e\��޷��瑮����E���m v'�z�?�,B��"r�j�U}�S"�4#��.�9�{�u]��|iA�/.	�z�U6J�N���o�� �dk�����;Hq/��oUL�α�E#��(KY:��V�;�s�"H���\��h
�w�����t��r�9����ļRc�fc��*.��ڌ�wY���o�1�/&�J���
�D3a�dH=�O�c7c�["6����
W��5��cD��[�]D�is���?3 ��чB=fz_�W4�������
�Fr�Go�A���]���A7��og���"�f!���Ġ��^	{M�n���O�n���Y��O.t���{��H�
�/�m��󪄴F��*��P��E
� G�#�zhPL,'�w��ثB�Z�ق�6��I��H�&��es݇��cUK��B�T9X���w�\p�A�V��V��1j�d`��˸����Ju`���uqj;p�ؽ<=�:��!�f�J�cСSéپ�m��ל0K럳�$F~Y������9�unѬ���#fqUT/-�oz��;ji�V�����2��}����]�C�ɰ�6�r8��Iդ��/�_d���A�=Ɗ}�ԑ2���d N+�
�r`�<w�(C���`��O�u<�Ѽ���6�	dڐHp�0#i����ZˇY6Y��at�(������i/H�"w�z�!����c�ӾiH>/v��8���Jgy�z�(u � �(�k.�8�]���Ou��������^��ܖ2�fiXHm�>�v�r��K�S�XS�+���R���o�I���'�o���@ ����$(���;)��!vMv�v���FiB$�C�s(z�.��ª���A����i<p���e�fC}"V�ts��gJ7}h~�;�|��
�,�p��IO>Y hw�%FX��P�t8J����zd��M,?�G�M6��e���H�U�5�o|��3��ޤ
���x�B��F;b�7<�2�+5y!���㭧�ůӊ�C�����
���XZ�}��狠�Ջ���i���Mm��.��e��G��/b�L�Ӥ����7��B�͢cy
��������U+Ǩ����|0���*�s%�Ee�/��i��R*!V���	�x�'C�7��M@T�0����~j�t��@�_s6|�7�7��B2�l�Oİ�쀎D=���k��yk��pr�<ڦ~���a;J��dZ��@,���*�c�c�F��t���e�Qd�ZQ4okz#KI�<���]�^O#��}�>L�$��=d��pz09D���3����J)3JJ�ȟ�����=��z������3Ƃ�m'b�Oh�Б�ɼ��S�y�$'������`A)>�*:^X����c�4��z�s���$j���q�yO�U32ۋT'�wy��7�{&�>��;罉U��Cm����x�ESS?"�~�&�O���6���4:�	�c
���(}����1 b|Fo�������]��W�����'�Z�>C����xm{FM��U��=�xw8��M��"�I�{V�B�8�s/�QQ��ӈ��[�]�Ѷ�b���2�e?��5m��!E`&$����*�VD�wB�tߥ� TSAN�ȴ��t6\�&�oS�����l�0'�ӿ7��2����A'�n=�h�ҷ����<5�6�\W��K��|"W�7Cn��}�b_�N"�w����q�2OT�c�>��IaD�1�|J�����/t��n�6c�p7խ�x�g���cP0��= B5*OI�"�K%E<�jߵ���Wv�&y�>r�%?�2�|�?����X��+�f��g ��!9K�k�.���x���W?sq�-}w,3C�F������ZB�`p(*��tz )�YV=Q�׻��^��ĵ��DU�=��'�Ym��A��'�#��n��C���R�����A��pr�����sT��!�H�}q�ɦ4��t�AYJM��p#�Ch�ޢ`B٥��+Zѳ-ik���Z黾?>V÷R�h�jՐ���j_!��|m�
D��޽�/��Wߐ�7 q��w�dj�9k�b4c���kW_oW�;�Xu�:�=PV+b8y�ی�u�25���5���߳�x+NC=��Lm���~�q����gu�<]'S`N"�r���3����n�:��/�EP8���N�J֖�]���fc��A�'g)�JktM�듙p�������,0�����ɐ���k�����	NB�rA���n��-<g�M�"��S��z�t�lL���P/G,�M7)�E=KT�yq]���f{u7�V�Ѫ��o.�����An���lMa̪�8e"�R��ZwF^�bė9p�p$�u��<���T�C�����Y34�z�t��|.�1�h��~\X�29am��Ş����R$h�2����Pk�x^5`�&utJ���Em�,�ôk�DsZZ1�d�}����h�u���Ǥ}����ܲ��j�oѮ�5�����/����"�VDG���V����r��ak1�B��߽��O��>fnwP�����6�r7�D����OH���44�:����d$6���.7a;�U��q���g�#�b]W�m>�>�d��TӜ忸/Z4���@C��'��Ƽ�����:��M�D����3R�����������=<���M88�b� ;:L�1ڠG>	��i#?��7@˅,�?�*�=���T(�6�AN����Z�tM�" ;���_a���`ڡq%���6���f��!9KQp�de&K���i�Ҁ V��_�lƑ����kEl�r��v����x��m�K��l	�)�AQn+ �͉��	��z�FP����?FP�5�_��ߊ :�x[7���	-�ζ������������>rܻ
�v��||��w������<����~O>!�]+t#�%ݙ�(�6Q�Jx������"%sdX��e�s��ݑ�q��ފ=��h�L;�4h{��\�ҒL��	�Ec??6��C�j���a��,L(�k��E�3v�Y2�] ��(3���#���G3�:��}C���E�z0�s�y�<�{G']rk����x�{����)|@eʔ6^{�Ǚ�X���nz�H���-�X�h�����Q��"����s��F��/��Ɉ48Ҝ��!1pv��O��;��f�q�P�%9 j2R� D�馏)���^}��ѡ�i������LR.a3 ��u�́�UI�Kq��:,?�@��������#C(��J�Q�=A��v��8���cŨ��l`�ǧ��X�������δ��#2��%����w��!�h��K5�L�g��T��@n�Ʃ�׌���.����x���yS��}B_�S��/�s/�Ic��jܒ	����w#��X`9UQ�
�
q'���R�F���xms����^�D��G�t�_��#�ƱX+X��Vp�nEkA�X[*��z�� ��@�-:�Chj��3=�.ac)�Vj�h� D~��q �g�)��"3z�Ѯq	H�\�=5�KV;�[*�:xv�!��R���e2�g0}�)���Y�śs�0"n6�
c,��AF��=������&�6Gy�h���_DP��ػn�$пa��@��w�	�;y��F;�5�wN0R�|���r%�k�=��
�B���/�w�Ac0�B��3��_l "%6��]U��:�N�]�jjq59-[�P]Pl+\�δ�r|
.zD��e���[(�����J�Ͼ�'�/`�.�O���7�@?��C�$WK�T�	$ٻ%�N	��*�){��Å��$������j� 9a�*�@p!I
Dd���d����3#��3���庺����QWw����D�K��Ǔ�|��dG��I��ial�x��`fs��^%� s�NV����T�3K]p�J���Gs��`ЧBYs��!���>7���)#U�Hr|��2���Y�RQ��0�/7���H��BKv�0�����Ĕ6܎�D����"�K��i2�o������N�
��*aM�ZE-g�h�U�|����� ;�ؑ���:���Z#?�_%�����j����[8��kY9�a���s���������L;�a�p9�}�f��H��A�+tme�ǰ��dL���ȋ��~�k"��q/�z!��9�$�N�D���f��a���afPcr��,Y��L�b�C%�"o۞�o��VN��-�*��M�G�t55�$�UF)pI`��1{�:f�Jj\��
�!M�.F`d�} �NՕc�!���������}��+��U6{��Rb��m�@Om����PL�^������s��S"�Ƃ>����*1/0|��"��݈~��ˀ����C3+�H_>��q�Ԗ���zc\�I���Ѕ���2>	�XhIm X@~s��X�1��p��gv��Yw_+��$)�J,S� \y��q���(�����?��|C�/��_p��(��� �ŎJ�cp��MBkH�~�q�K��K��{
�Ģ}|rHl��&� �@�U���	=��7	-� �l�ν��"vr�0A�z�S��m�p&u}eE�����7k`�����=#��@���։sV9����,���Hy� ��/-��M���d}��e�
(�����ZQp�S�(���\�2�!�t*�,s�x}��K�7�[Y5owY��ҰN���-� �a[���'$���S��e"���.{��>	*F�(��7+SŹ�����JY�n��(�L:�H{�Q�((vi%W�	K<6z�L�����h��Y.]"�:In��	!�ƨ��-���v�ˑx\�	A~��)��!e�\4<0�����L/��iD�~Z)��{�����n������� ������.:������n�(6)@�钭������[`�)W���t���)���f�4���oN����4��r���хH�j�ڪ2���1(:�rw	��k3�1�mLƝP�p�r������[J�@��8`1l��7��怪k�ڪ���g�>O�?W�\I���v�M��p�|�-6��đ[U�ә���yÉA^ˬp����_6O]�l[q�t�]���q�r�um�fx!ӊ&���{p�VK��+�y)�Q��y�ǚl���HHK�nQ�G}|Vu������G$��!�o��.{�����q+\��(~XS%�k���r-\Hf�w=a�6Xp���f����ѧ�>�h�w�Y��~�75D�QR�;ُj�����Ck�L�-��@�&Ms*���Щ��1�n7v���8u�7��	�[f^)XA<��#�sw~�����*�
7���{b q#��MP�9�}�,`&bs^��%%0B/�;_W�#8�&a_z̨x�lA.<�NnsSy�$�S#͝�T-�ֹ2B���6F�I l#)�^��U�K����~�&��,��a�2�6�@J�j�M6^��z�	Ń�����H��.P��KQ ��l��)ɺm��ϊ�7���F�d��Zm��*���6�E�~c���w\�T���<]���T���'f��d���W�M'*3c�z�m �B�"X}�S�hʫo�%]F�M��E�I�]X�g@��	gv���S�r��@ŀE��?�5�q���Q����y�@A�{̹��y/�|ѫ������׀���Sg�{��Z����.�,γ��GmŸ�WFħ����f�@
V�������n�����n3���1�ڕ���]�}^8� �NM�
 1aX&�?����%mt/b{��y�G�]K��:1�4FJ�߅�y��5���L��Z]��V
�3�"|y薵���Vt�wT{�;c�������^�8��6���Z1�4D�"���Z)|��:P����oz!�Ն��Ș�b�/;_ �|\j����Q���E�c�Q�U�f��҂2?~�!S[�)#�c�)pI45l��q&��J�E��_8u��3�	p{!}vAIHNS�ا���z w�/�}L�lPă=��G��n�>��jw�~Yht�/���!�
R����V�V�K����.���y�`�0�1��Ӡҫ�	�>����bi΃�G�7%���B���Ɩ���Mb3������oP֛�vCY�xW4������uhңӢnV�o�<T�R�%U��^+1ujjº�g!x	J���PU
��0=*Tq��8=Ċ'»l�f���ť�����ܤ�����}�C*\�t�����R�#U������H�&�2��e��\��ҎoӬ�Xb���8'5���' S�jdاVl������,FgI���,�!����j[G��ֆ�13ΔA���
���p=�T��g?�TPl!��H%�65,�t-�����m���D����-����ݭ�6U /��q��wy�,����lڤ��wռ�72���Bj�%[
�!J<f�C���\炲a_x�X����j�sBU�If�Ň6�)����5�|W-᥾O�h�x�7�sb�6+gܛt���,�U��|Na���L��,@L�)[��%-(\�e�'�g͎�@�4��_]�����ݗsPǤ�7�2b5���-5���BE�n־��J�^��׾�,����)}�̇����U�e��H��6ߑ1C&�a�e`4�8s(�Lp$h�E�_�T�����n}^>4U�3&7~L�Q���(�us���tՇ۝/������n��1ϒ��w�
y�G��:�@E�I�/�G��Dr�q��%м�/��A� A�h�y���������3�ոo��*�|�%����S6F��Tb��c  ��ki|^-�d�
&���pj�"*�[���
B��<g�)���.U�q������V��z(U�<������qV�U�@DB���e��5��TE��F6��ˎ�Y���b����g�ExM�9���Y�I-���U�J3�D:-9 A�e�^+B@T:N��F?�ڱXZ���jZV���}��ݢڳ1&���Uc�7��wa�L���Ȁ����඀��9�h�JE���@�\^��ɦ����[����Óy8��g�"uxӾ����L�����k�UU�n2yz����������@���5�:5`[�%�$Qa�@����+J41J5��N�,��Mj�i����|x�/a�ש��H�{�����q�z
O�}Dh�H4b[1l����O�g��@7g��������6���l ��n ���?z�ݗ�Q����SPK�P^�
�ShH�0Bc&[�vG.`kL�썑l$5���]P�e�2l���F�@S:>n���ɣ(ǟ{4C�A�U 7o��O�)M(o�A�v�-�)��y��D�4=%���(���_��?R�a�\<�����*M��o�[{a|�.E�����Ia��4n����j���.^P��ߓ�~i+D���C,�;�&Q4�"�.us���d=�8���B{������1�u6�tt��ނ9�	��Tפ�<K���2b�9A�W�L~xx�K�"M� -�N5�A�n��_��N9��[ ���Od�A��Q�6��:�}U2q��$q��_�� (��|u����Ŋ�w�>���A��U��0gXJ�l^W�`+W�jx;v;S�Eޜ(�,ª��'PQ��F�~�$qyBw\>Y⫇�XP�T9?�o�F�%v<�$�V.ŷ��ޟov�>��삐p.���M����k�����
���˙�n�ӓ3��j/���1�+0J�fP�j���|HՉ�-@n�2����3�qŢ�d�%fU#��;S�������<	۰�Q{^t���a�Uxi��� ��3�p6d�>�	^�!�aPT����b�\'��m���N-���kY�c<[���]\�� ���׌At1h�0��}/m�������J&VTe"��@��G�ş�$��pTފ@�P�M �隃{n�[�o�8�/�&��09����SA���z,�S=ֶ2����e��Cc϶�[��EGh�_liK��P�_J�Eu�gx�B�<QM�raX���UJ�����D,+���e��5��L8�G~U:j8��Q�+����\�*���I[��j7����pT(�ܲ�
��f�������W�{U*}jc���A����4��M�@�5]��Z��?Y��2��}���}*�������[�j��>� ��S����j�SP,���0�¶_�(�Cq\���d���>pxR�Me�sy�tUK���ޥ��ܨфQ���t��F$_/�S2`��ܧ`�O=ֺ�f�T��O����wGn)c��Q��a����zE���fg����6R'N�!8%px��g�?I�VL���p�"���>QO��U�%����~X��r���+c���2���n�8�=-�mJ.�=p��4J�����w�p��O��3����8�4���`���6{`@GX�~(�1'mI� |Zj2m����=�Yn��ϣ�a�k��&�,�-f��H��i-1�y}v"�8h�b"k�V��E���k�cݕ �gE�����W�-���������wt�i�ڐ�pF⃈'��3��n'}��q���B=]}���v�a/x��f;e��}Ų�g��+7��cr<h�N��s�G�<�q���g����tK��Vc��0���ZunT��?�o-A������:��4��ɐ��v��@�=O��IVQ�y� �,�p\��{xy�x�����%�����B����Xѝ/O�O�+){8�K�|����?:��;�[��l\b����u��H"u�E����+mO�4oN�9ԗ��ķ� z�Q���fy�e� ��-N�dO
�"8��7$��4�<�i�Z�7�b�243�:=U��]����2�z�7�42�]��S�g>c���9�����X��%_͋��2i͛-"����5���}|��]�ۥ[UXJ��`G�u_<+Fs�����[(�v������(�$��X1�wU�������[��������5	`�.\a�����hf�>>�PNR~�\�{��$�C6S +U����$���f�4��N�������w1WeMT/�}t�u�T�F���@���q�	�H�>�n�C�rd3G�(؄Jp""yD���Z�)�fA�f˹�d$4�Kr;��NW�9�m,�:&M��]a���C��et��ICw*jR�����#1\��?����^���n�L��Ϥ�K)�n�Qy��Sz�ScX�+��-��|�[0��ዌ����Q�L?vГJ�x:�~�OF`�ݑy���v�^�w�3{f/�j����ȗğa�.���74q�hRŘ[�^(Q^����L�[���^Az�R�F �2��>��iX7b}�]��-�~C����a�[�����S|�V&�0�g�;դ�.�]��r�l��ٶVDd/�����Q��v�GOȷ����N-�΁�H�(�*��|ʫk���e�9al3��WQ9�/���^����"u�
�F��������kl������wGQ����i��LGK��z����
'��g,w3������J�t�7����_Ch�P��q� WF����w�( �F{ ���7�����q�U�ԧ���C���0�`��x�,n�r���q+fgT{H �|:O�?�ع��t�L}�pHh)����[�F�	�>*`<:#8*~`g�#����3�'���9�b��{b<E��`�D��7eڷU�]6�M*�*��H�:���u;Vw]��3�Ԉ��Z&�c$Hr4��cL�]��I�?\��~?�7! ��f�Y'���$���^�n�W� �0�`�8�K��Q�ǧ������ �\=q��V�n��
�O;c��^�(��K��O#8���oۆ��l�A�|�Pޠ�TK�h>[4<����je��"����7�\�Ir�>��}8�HM���DmGvot|4N�NK]L��
 G�e]~=ܡޣ$t(�\�tJ�ԇ���`_F�T�٣�6Y�x�����8�J�߼����8��kC�j�מ�g|;�OLl��	e�m��-��z�6�f���;�r��v��&Q�Y���5{DS��7�Պ�����c
b��F*I����6�bG3,	 <�'��Q�Yf�L�������@��;�2�d��v^p�Ă+ �X8���3f����_�^��k����`'���=��=���Y����W��_�3ۥ�O�B�&�$�*X�,��/=,�\5����^F�R����X�rx�j��J��LY�2�����Bpu�er!��+MS��O"�}v��Z�P7z�a\�X���D�]U���X��F�����}�B�s'���3]��r�;d���<�����컬b׹z�&�u;4��͐�'D^+S'���rc���=9i�x���澸a�G��j��*_��b�7ds��cI�r��lfa��FK��6갬obصl�9A�Y�U%
��;�&�U3%��M[�憮>c X]0��W�aՃ95`�1E��ϳ7	ʏpU�-���3�����;��~��a%@��$�M�p9�XO��)0����G;L���J9�
�g�2W{�p~�~F����l�7�i��8���Ն:Gjҡ�E���?�5���ܤ;�_Th���Fk�s�ԾTB)e{���Y�w�ث�A��M�pm�Q抩\�z(.��6?��>�4��j�n��cM�� $dc�b"2ż��o�X=��g\5����H���юj�|�o�>���Ĭ��!i���|�s��0����I��g�F��L�۸�D<xmmp�߰a�o��F���4�P��5(� srS⫦)CT��y��󒙦�`�@}#M��s�PԠ�� ��⻹+��8�t:�B��	[�@G���]���ó�ufIM��Td�l:�nE;U��{CUxK��/>w�i��PZ��ȡ��z�BF�S"SKL�b���bo?<��猑�0M[$@_�:��8ડ=qH�U�`�hтU)2h�!�%%@3����W��9kv�4g�B�T��~{�N�Z�o���RX}֏���S;�����q�`@cD<f���2�ЁF|�b<�l���1����a��:$�{��f�-����ف�F��YS@;/��q7��Pv��x~c��xő �r7P����e����CI^���yK�~Q��,���V��FJ3�9G�EZ������}?c�,�6��UM[�����zs>>�2���sC�되&�O(�1�G��#��w!jv�Y	�'!Ƞ1����;�g���Ϳ^��b�g�#>�E�v��=J�_5[�m�I~�].����,*CɋP��W�}vV��F�#��r�B�wMe$BXu��3��`�����X	�=��qF�2��BZʄ՗4���Y��;��3XV�qg�m��m�mb�j'dw�Ӯ^����ɣ�C�O��~���P��=a�Im��0 �vf;D32S#)��Ll�QQL�/Q��(F2w3U���N��m����QE�x��%W��F)=��H ��	ҁ+�Y�@��p�5K3�|v�C�H�ڿ�Wb��[�Y�q���_��`�Md!�-h��kU�l?k1�R5�
��@����:�f֝KXA[�78�)�]L����2�퀛V[�iq|xg��ɋ�Wr���e��D��ᄆid&Y1���s%��ه�4*z�J�2���~���s[�b�g�E͉{����0���n:*0�Ğ��������Wr5��&H�u�'l��+n�P���*�2<�F�Lٙ��7+�%��<ˉ|��9�J���n�L�K����U�x�C����%{duХ�ʼ�ٔq<r�y̻����k!t�HjG�x��Ŵr^z-[�;�;B�k���&h��p+�_ȯ>ô/��,�|p���pЫ����6`_P�]�<, ��ҷ%���$ˊr�K��Z��@������;#���$��k�G��D8�/��Ҏ"w #��9�;���~�}�^���Bw�`�A��,�����X�7"L��m���e��^�e�q��|! �ͧ7�#�l�0�_�m�%#2�jz�?��7@��uȤr���pƟW��� ���O�T�s^J���$�UU�R{���]��P��qjyú�o�cT��%Z�Q�`�.B�0�'.Y���'�%S,��3.�a�������{�7�
��^��<�,:[���_uEK��ޘ#;w�ϴ��pև-;g���<;�cط�٥K����"��[)�L��l���[\S�0��E1tk7��_�6-����������ey���9!���~�猾T�!�	�B�R�Ṅ���>��m����`�4��S��#�{����#}���,B)�M9�E��.q�4�bΥn��ᙳ��,�i�q�x}���Y��zu���48��P�{F�qsj����US^l+[A�pK$}ޖ��wgҏ3˺��b/�aW2t��P��2��)'���Z��Z�*716�h4ei���y]�F��wt�OF2�bw��Nd	��'Q����(2�:㧕��淯��+ָ"[�s��J�b�����.�*���!� >�uU'ΡJ�����*�K�k}T�S`�f�ݹH�h�6��0'�\0��}�p��=�I%�^K��	A3�G1;�[���]�[�/u�$�O &�A�;L�t˶1^�8��
�|&5\Ǜ���ވi%8*P�.�F3���p7n]��Z�\����PE&RgKd|א;����T��wu�7X�����;����E��W%�^Wٛ�lx��]�an��Ji}��;FSCIJp~Q�%4�1�%��0����q�E-	�ȸ��v-5
)}�L:���.f�-�!��E�!�cz �򡭤�lN1�ԥ�O]T9+��z�~S���ÊN��#�_I����]bx?����U����qE\�7峮g�l��)VQv�1қj��Ӯ9��ifk�XBՅA���4�� "
]��}`�	L��r�//����3D�D�U��@0yU����#���(�W���ڀ�ۂ��� �$S��\.���m/(��$5��vd��o�k�np���H	pG��0��|Q}�����zJ	z�<?�-φ��߂�O��B�	��r��>:zk<zvv��s3zP"bk|���+os}XeMF�H
�V�o�f�G�kY�kω��(]����?T��ޣ��U�o&�ԉ�������]o�|F���j$Fl�ܭ�=4Y�x���=�:%Z<��c��}Q��Fgp�T5�� �]�%���z��K�{z�̱[���Z�$�z#Y�n�j�R[�^-�-��H�4I�+Ծ]�n��%ꚳ����f$�A���su�)�����w�ip���~�ku�1.<�f�>��/�Ӭ�����˖q|%ɏ{�J��������%�]� �'�r�D��^I��~#jM�t_@�h�r]6����'��<���d]E��� VQ}M�|��RL���ʉ�)&�Ac2b�k \'����R���E�-ݖ�&{��(c.?[m��Ť�P`o��������kr�� �] 3����B��wu��}���%����hcx1��TS���kH̀iG�m�>��K��f�i����z}�}�zYz���������UT���M`��Dם��)���L�����'!HH�(�~Jy�Wi,�P9\���2�SD�1JlGu@0�ɶZF��	5kl���Ԧ��+�4�/��U��o���rH�kbP����ٻ�T�!����)eB��p?2nL���-�0�	�<_͕r�'I���&$Ut�l��u�`��唃Q�V0��e���k���mI/5tӺӿ��� "Vy�j�K�84/�E���B��_�}�L~h\QC����R�L7b�	�Y3����%������X�e��K����x?�vof�~4�w���|��jT*^����V�j�Qm�hg���wpH:�\/%�q�VH�y�Qh�`&0Hޘ�szF�U�6�*���w�[V�XB���n�:��L8�W:ϠU"�\�-c�^��`q,�0�`������פI�-�f���~�o�!�\!'��rnu�ei�	��w��}(�h ����2q=��
F�i�e5�%�������S��S���Zp�9"�u�|\�� ��@0s\a�`bIC:6˃�1d!�<�lq)D*qm�h�S�~�=w���2�,��Z����0��y�/�R�A9[R6����[����r�����n[�Ņ5��"�#��/�AQy�:t�L�E�l�����rP��[Ȁ@ k�pՕ��?B��`��s���6`���oR!2�����F͂�-�N2`�{CN�G��.s�G�<�O��ɖ �-xJ'�%��f�.������:�E��t�]o/�\}p)NI���ғ�\��a{n"szP�:Q�&�a.��h"���y��qW�z�k�p�>��z��nc��s��$�:!�>խ�wv��X�6���V�<+��B�O}�, ���s	Q��a9�!sMl*�Ɨ�"M�ֹl�υP�8�LON� ^g�����Xi;M�9� #��b*<�Ɠ� �� �/��z,���,��bO���8=B�BV�7��m3�)��]z1r����'Ӿ����v������/���J�.í7SJ�X�0G�K�%Li�sfD�'��8��i�(��ż��a�a�o6c�+2Jr�>���Jt���<VB�������מ%6��V6��S9���'���5�ڣ$]e(�*^ ���x�,��!�gD�(�ye�.8��m�������z���9ɯ�a���M�~������O���"�[N5��/�zvj�ivjѪy	�����Z*�[������o[�g��/����US�ƣV�Ӏf
?��RR��]�pu���Xǌ�wTӅ~DAp(�T�l���� u�w|B�����~2�_k���| -��&���oP^����C��vM���˟�@�k.��e�y��� |Р�lTr'�@_��V�3Y�1���J_���U�] �4�d��=�b��݆���Z�劲�;:���;(5'����M�x7�d:�	����[�s�
>��m�"�-��:0�M�G#Y#�R�ȳ
���sǹ�B��.9C\w�Z��L���
V�u�&X~�? ��	Zs��u��Y�6�	N���8��e���;l�ཙ�%�Q���9�Վ�a�`��YK�.��f�������Q����>GZ�X��c� �Z�b�v�9�������[��LPM?3
�\�a�מ�&�p�lN��'���R�*�I@Ob,s)�4NK�
�3.�2����C�{�d�f�mB�k���$�����<��Wz!�RX�e���+�?&m��}����a��8����&G��z�W�����q	+<G�yb�(01B����nq������C��F$h!_���r�H��hQ�T�uh��҃�9Ϧ�a���p�G�6|I�� ��O�� rhk�!�:�����Ǯ`�M��2HI�H{ʓ����0���<�V80��H�'$<[���(��	�aN56��3�C���/�9h��d����J���c�#�	^F9ﺖ������O��z2�m���ڱ80,p2��P���bf��;W�U��i9¨z!�R� ������h�롬���3�՜��(,��,|
�mv��˗�.;^]ܹb�8��((���I5F�cX�d��y&�4�tk&��<p���G�u1�3C�ޅ�L�JTd7����;'�P!S�6�²]/3��,VW���@ZI	��������$ZCa�������	Y	PǓO�hTNM̌��į�Q��;Ɓ����o���u9��n
j�51��>�XY8s`%Ƕ[=���0ߔ�-�:5o��Ix���]�-v��qk�c�f��a/C�@?M0��] N��o��t�uZ<���u�g��DA�8ەa�uzC��<3;�����_�z�����	�V�0���[$׽�sט�<'�ez���}�$h	�'�m�^�'B`�m���`$�䀉k'E�2Es��TN�!R�z~��h=!F����-�@���?r��z����Á�T��-VL5��]��i�n3f�Q�p�9N��ȥnW2��5�х\���d�?�s��[� ����$��RM�����`��k�'Z�s㹏��c�� �ڵ�� ��"�J󇜪o2���7>SbA"�v�+����� �"]�5�/����[+w/4%�zc���S�9�Y	���W3̆�w�HpmR-�1kpv�GN�q��#с?�M�W���"{�D���nh7I	��Yo�{�1��/�ަ���Ѳ�j��dʓ����ϞxY��L΍Ihh�Ӏ(�[�WB ��Cf�����3Щ)�H�<�S9F���Q*R���igP:��@_ :�c�0��+�b�6��>�,��ߧ�|4�ɵ:;�Ur�R�痒m�z�L�>s�#�_C��3ى?��^�eDz�o�g�\X��P��Ǥ�QD۸�K��*Tg�ʎe��<a��	���gt��K+�C�kzj��LJ����4���`��f`=���/~�_�hIC�gDpV�꽹�9Z�~rG�T���=��v�2��@}s�_9,