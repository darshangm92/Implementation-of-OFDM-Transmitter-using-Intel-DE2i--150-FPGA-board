��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J7���zZ�3������B��h�Y!,�c�k������o�!sz>i��(l�N�b�.��t�X��PƉ��"_��b��O��VdnH���4S��ޟ��'�S1<�@�m���?�#�FZF|�8�G�w���>���Ï{2�<�k�@YBZ����ϩp⾕R�UB�!;U2��O�K��f��^M��J,��3����j3* ?}{��1�
�c*���`�������+k���e��/?˰��%8�W�L��)�[C���=R�;R���8L�0�^�����B�+�c���j�:��h)�g�xQM0g
xE`���Y��Q7�vO���9<��Fc�R�\���`O}�}ĕ��
��jR�)y_%�+�]�b�k7�[ټ��KLz�?BY��7d�t���Uu���F��p7��^+p����n����@_�k&8�櫣=�<�h�g�Щ%٤�B%��/�b�'��t��r�I}N�G|���o��i�j�7لY1�|ߠD�~7.b��z�3����(b��BuU����/s���c��KEM���%��[�:���6Q��T|�}695�~�x�Bj�]�j 	V�MH���+�l��j]>�ѴF�ר�bLV��B����k\
C5�N��k���b�S�!�f'=�[��utr� �1���I�a��c� �ty��W~�"�B��q/X#���\���.��%�hּ�Y��> >�.Bv��wimHC�U�ٙ:�h>_%=��au�`B�or(��_!=�TE�Y"ٸb��+�Tu�#��=ӣ���F�}���@�aTɪ;�6=-���~�7�� �bɇ��\X�����)��i`�E�(�e"Ҁ�UG'�N�	����T�ձ*�|��k���@Z�����^<�	����u@Y��pI�� ��x�(�n�mݹ&.:����a�P���(��s�"�>�15#E9oo�����ur�(x���0�B����T�OOnr���.�1�IQ���i�
iF(�$넣 ����އm�&��l�$�J�9�4O�}����Ӷ�c���� �� �;�	�����&cI��m�fx�FZ:���7���1��;�N��[���rB�t������=�73�����76�T�2�3��y=�$��f3�����U�*�đ��[�+���3{�������D���w+�<���\�K���*(�t˚�]0�3�ǩ��pb SN�E � a	^�5��4�
�eft4IW0:�-s��0d_^��m���,k��د�%�ip4�}�n���W	�����hv� $��U,1� zl�^����NtF4%����h�;�r��G�}���^x*��Rq��j|!����>2��k�=�7�Z�3�B�j�kL��Ǚ�%�n�z��bR_�r�柏���g:P����q���?1Y�>W����3�P�S�R)P��1��98z���b�{cY�"�����Ij���o�����Hݳ����RR�m�cے�:����	=��摻W��@�σ��⻞#Ȯ�	v�w�hyE�i��@x�.r?)�j�<���PE[4��E������E�u��S塒vS����G�3�pѷ�QI�by�!��+��;������+���"��3��K��ѦHB�p�|7u,\���U_%��e��e�,C��5^`jR�?���Wlɭ���qI�J�ݡ�a�*y�HﱢB�|��.��%Z��2v�bT��I�\���ͅf�w�~%^J��[�Ux��3v7J[�a����d�ؘ+�P���xʊ1	h�~>wMn.�p)���L)�|	�40����!���,;a\�ĺ�P:�������A?��DJ�Z:uE4F-@;�P=�{��Uvm�jg޵�^y�!��*��d.\Ko^�~�3���O�~@�z�#�(6O?wnB��)�e��iqm�wN��߮�eJf�$���b�!Ho��m0|�F�����e�K\�����!�*���ї��t����.WbS��}��j�5�n^�WlkF�Y#���� (ng&st���sk.L��٘��jf%�Qr���e����ؖ�շ=w1^(�K�>Y��'C������k�a���xR��+W���P;�)�����0��GÅ���Q���)�[�e%̵!�Sl}�Aԝ�B6R:6@�c�(�8�U~��L�����tR��5�Tz�|T� �yJ�<�T*�_T❞��QZ��9����]��
��p:h��Ӷ��{s|/o�Y�k�[�P�?�#�ν�z�0��ͮ*�GfH(I��CZȅ�C5Ջc�ɬ����F6���s�ߧ���~U	�1F�e=�3��)�n�w�D�W6I�����ew��]Xi=�����L���y�2����Z5];:�Fʅ��'#QT�l8T�ՊI�U�w����b�PL�����ZP)��{3����wG�"'A��a��k�h6B �^Y\aw��-�u�����
� ��w���/z��3�U|'�%�w��QF��ݙ0�\k��!lOf/��������iL��:3�|e�ւ 5�A�h��u(�/��5EE���B��5\�q��l(�%;4O�!8�i��]��������׏�=6�FSQ���>"}�\{���롽���h�JI�q�/�-JTk��:�Zt���L��Fw�_���g�t}��� ��e&#<Ce�4�U	8��-��%�%��f�s]�o�o�����?�Bk9�o�O0�ņx2۔T��ҍ���L�.�j��Y򹚙{!�vb`Z�D���r��p�=#6x��Kz;��紵%�2�9������_&ؐ��Bv%���
�M��+9p�6��9�
���v�d3&=,6��&ߪ����%N��=��ǝ�3�T����%n��Q°?�|!�=@�7m.[�\�h}s�;¾���6m��2���B�8�QRMhs�7��h�}��:#a��OQ������gT��O���z�Ɏ�O"��a���"K�ub�_�΃Y�4�Q�ŃC�3�h���Vx?S񃹵9�n�S��<��P�,b�6��� ~�(�E��-0���=��p�$�L�����E� �;L8�q��t���>�-���)Yr!Ӟ���v]Z�䲙0�+-�1R[wm[;8���T�N�Im(�(���cƼ������e�+� �"��=�5�] ql�'�i�j��lF� ҿ�y�<ugf��n◀'0�Ș6����8������8�vD�
w�'q�{�9�M�,���T'��7j�Ù�@a��q:^���Ѫ�(��F�&A��qz����i"�%4��<�=��7��Δ�oo�"D@~��^�J���Ź�z��ѼRj�J����=}�����T�H2b�y�#EЂ	��������u����4܀��z2 �7�~T���/�O3�r_�R���im�_<�<Vs�Kp"��K �-q��iz�����zPDT��������`J��8k��/��Ißڥ��CH�����u�~��?��h��R��с #/Ȁ��7Ï�/��7�R��D��	����e+���k}7=a*�H��ӳ�%��*7����)��9���Ϥ\;}����."@Mعm�r�:�Ű�Yo13x�������D]�-*�y���N���{A��&^��T�8D�q�+3��1���Oj��}��S����4ƛ Q� ҋ�q�Y]�QFF�8	�`j���C
�˵��e��^��M�]��K�ȼD�/���o��ƻZ<�-q�n^/�m�s����n���b�KrV��gAH:��pr�j��f��9�&\q
�7���	J����4�����^��iu#a9���HI{a,,#^���`&@.%q���R�I��Iі6"/Aܵ99�J�[j��GkR�v�W�	%Dr
k��� ��Q���y66����Ы�}��Hg�WN2X�b�p<H����Q��D�z��F
���A2���=x^ݱ
^}Ғ���s- 8)���%�])�_(� qx@�m6d������]D�g�9�u*���:!�W�?B���,�A>�O�Du���ؘ"��m:�2�\<��/K�Z82\,j�b��-����e)��;#�/�������3#��7�|���͘Tµ���v��92[���g0��"!�xmzS�0+#x�/��|�i�} R:�dUR����y]f.�1zi�4�h��JBt��A��Z�ĨK��o �;- 2ũ�`�' �~�3�L
����Œ�L��ߘ�kJ)�Z�$�<�Y�f)rj�Y~B�	Yc� �o�
�~e��?�"a�$��w/)����/Yɓ3�l9������y|n��7�o��o8O��@חڬ�����BXҾ���7J�ڰ����^�%���28��1�4m6^��������'z��5�A��^�L[��1�kX��>1m� ��5G*�w�+���!�EC�@�LR�ć�_��S)�!�_!E�����7���ug3�����Ҥ��'�|�U�9��S�w~{r�	z4��gw�����\�8x\UL�ކ����BfB2�2+�Eo����a]���(���@o��)�Yf�c�ˈ&1�	�xxUA�k�����H>i9��g��؝² -r�����"�i���]��;:a��)c�[��^�%t-��i�3j��x��(�PI+d�^ί�v��ݼ���V��q��{�c���:}� �D����WP�˯*+�j�9�;߃�w
��aȑ��v<zOp�h�ce--j��I�0�^e�K���`�W�`����ӨyNZER���q�C����]��ˑGɠ��1/`,d� [�;u�T���5'��`?e�՜#&rS�z�����K���c��� vl6���8�Q�4�k�6���_f�#%�َ:�U�6��x����Dz���@ۼ�H8�e���^��j}�F�c�w}�4%��EJ��T��9G
�'M���s��
��Kl�b Q^��;m"^��rJ��4���Φs��O=|����_�%�������@�}��i���:?�à��'-��ҧ��#;�8~C��撇����5-|&K-���[��؂�f��M��ZM�M�
�&��T����rj<�5�\���Q�{�F�v��$���Զ$�-�|Ŕ%&�ᗝ����R�nX��t'+B�Y��&�{5��E��vah[~���PR��3;Υ���	�0��2���1 R�oɆj��x%�[�L�g�9���W@:iC���Cm4K���g$Y���-�\V.N��o����!5t/��_͡<s�#ѵ3l0M�М1()U>��屻^���iN���B�:u����ǰ���V8�W����������yFP�O��~\)�oS
ha�w6!jX~.��������&U�C�� ���Sso�H=�E��䋖�_�m����� Y�DHC�<�[7���֎�j��(�h")�I<�	4Ec8����*D�Y���i�l�&��\��kL\�'t� �D/=;��9��T�����zt����EN���܂8���ޛ�׉P�Y���5��%���
� S	����ju�V��g!�hy�ab�W�~ּ����e/"!4Je-�)�
���{��b�s�{����n��Xp���&1��يj2�R�
M����4�:2ơ��dXF�VG	3,�v�mWx���eՃ������P�x����B�f��T��b;�W� ��MK&�~L]��V���R�9�M�V㑄�8siz�h���5�^�h*;�{x�d�>6����@/�IR�B�*x#�&w�/(��6pR�u>���dx�7-�2,���=s���D�`�B��Q����	�UN,�3��!��s#���%��Y���G��k
������oҳ�Z��/��i^m��HXȏ�5�����g6�d��Y��)ne��2޿^�0����_Ĉ,~V��^��S����L��q/���Y���e��	l�� ��o���1��Z��n���[��$������]�/�H��u]A6��Ɏ�|6 V�$8�`J!�1S��Uʇ��Ĭ�q�;�(۝�P���}f���K)`jL�.fnX�ę�&�6�3.�7�������.)����}�KUB������nXm ��o�Ze��IqlV�d�� S�jρ�*j��=����7�賩�D��Ϛ�xO9�8��$֢���+�K�N���h�)9c914�yv��JܗJS~R���� <��y$��ήX��>�.�T�CvMMQ;|ל�h��	"A�X\9h�<W��t�VW*[\\V@%};�Q�
�	�뒠`Q�aD_vßS�x(cw��Vi�(%
������R�,��^C����6GsÙŵ0JpF&�=�'RrL��e�w@J��2zI3R���$R;_����-�4p�'D㹴�-=Ḏf�]�9�7h�v�hp�����whk2E�<���yt1S��ַ��K٠�^�L��y�Ӄ������yfN��������5v�:���s�/��{�k�u�7ɝ��ѷK�'
g�d>�����ٷ*�/��P�����/7r��H�&[H��G�y�P��Z�:;�'7*��fm��|b�%u�C\L@:�G�3s����H_0+v��:hD��l1a��:a	'�WTB�P�Qt�����7g\Z����q-��>��ѻ0�>e;��A3j
�QBNu@��;�~��߃Ԡ;''���;ˏ��z���آ���*�E�14�'���*Y<�)NX�>(m����/Gw*��Y6�
����ȓ�L�0<���GP������ڳ'��ʤ ����fi�����!�{� ,}�O}PH�cs�����aXd��C�UG��Ƒb���>b ����eq�����PC3���6�B9m���КY�Ǌ뀃MF�=p$d`5�y��e�!�hE�?�{��<�h�M����:�����r����ab!Y;�%���^9G�=$W'5�0�R���w��e>�'v�2o��C5?�B����Vh�ߐ]�|	�u����%�%iOK��5�Ƙ N���I#��G��� ���aE3p5�ю4�S�~	��[@������3����p^Ř��Lʰ-*���v>r��3��P�5�V�	�W"�4gN�~�OS�ư��rI�h�/?G$?�ݮ�H,V1y_�t�8�Q�I{�jR���1T�|(���3AךI��vA�C�� �9d�l����6�~�����\e}�(T�xQ�x���YJ���D�gċ-�'�E�&�sh�m[�"f���XG�\��`��(��!?v�Y%�wz�͇��Q�8�AY-�x����_K�Y�WE����JU���B4�Zw�4�Pq�J1-	]5��m��k���FZ��4'Jǔ��jng��p����C"��adw/�����%�k��OG���,�[���n0;,��$����,5�{�rb�\�����-cv����ݲr6@�$:�_>���J�,���|P80�ltiS��N��Rp(ȫ���"�c�a"%�E'����}(����q���m�L����v��f��Z�1J�n��d6q�a�`�쵅S��$wU�ղR�|zk��r/	��<�����"��e�'�Q���ue�j�}\�JP���n�UbiS*��0
��Etc���|�+@[m��d�rܮv�p�/x��T�DWZO��2:Q��Kw�w�pp��J���]C�q�`�"Ϣ��a��N�":�%�f�7^�O�ΛU�n�^2�4��ho�p@)���3��i�
��Xq�ʜx5/�%�FA�,0��+�fw9�&Q�83�=/�8��lu�� �|��:�*�o��F�����B@FD��w�"�)޼�����=@��q.�ƕ�hit���
�L#m��fo�fyx�z�|�Nne
���w��s)u`C+<_���=��M�L��?^�N����w�"cMFX�ˋj*�C&�CH4fõ��g8*�d���U�R4uI�j��i���-?~X�4Ez����+�[�"Y��ӷ�`]���&�č��l��?�Ts��uryWv��$�%��:�PcJ� �;�<w����j0��2w\h�}�H��T�g��k-S�B�����lr$t�ϕd�ʝJ�� ���D�k�%@�;6*�=�� �ӥ�>H���w8�^^^�;97�����u�&T���`<E~E�J�<��PS�����_��cZ���ؕ�b� ��IxH����	�w���2�F��Ib@x�����d���
�)xa�h1l���Q�ï|�iG��ʌi1e�AkӁ�ǐx�Ǎ=R�@[��l�5��7Mw�ڡr�n]�Њ�y��d�!�n�(67dwM��~�P��-�$g��n'lt,�a���+I&~)�Y���kH�<V�)�3�"��2-��Qvoc���V.#%[^-2��7�~���\���:1�x[�/�T�n2ea���S@f%�`��@�N�Gg�0u�w�6Q�w�2D����l,U퍬��'�yL,$�3#L�Y]]�W�9I�܉�M��Q%�!7�Xv�:�'>�խk�R�0*`����s�T�#���\z��3������B��qT�S�
�-1��������\t����阇�%q� �D�q��� �J[�j�g_)h".&&\.%�1�(M�����F��a�:�Z�،혻����k8,��zƍ�	�e�i��H� fӔ-���_�e�wǌD�<�SC���0!l�X��%�\�_g�nQ8��U'u���b��{4s�&Rm[/
�p`~�Ȱ��^9��v�����iM��tBǉ��V%�2�!IS����M���/g&>�R�����xVKܧ�6Y��a��@�{R6�������V$b�h����6aTC��J�����jL�P_�Q�d�d�j�3�%#���7���%���-��g�ky��Y6ǭ���E��e�A �Ĵ�숮j-��(s<�"$'��f�kpPr�٪�t[���;QK����Y$w���qh����U"L�sr$kdK�� �|(g��9��z��~wn	d��C������=l�4�kz�,���WE;E���P���s�K�,������Dw�PH������9�طp	VũI'"l�"�h6%
{���������a-���M����$��n=r�S~_H./���ᬖ���"�9�a/3�1ͻ[�����e�C@��Ջ�]�5`wY��Q��KR,���V��$���C;����������.�QK�|9��[hBk�6���]R�,H�4������ ��oh/�7��4�i�ns�/� s���xy�&����Ү��W�SO��:_L���K��L�Y�S��u��@Q�<s?5��
��ǅ������eK�+��j�r�4n +���#;����D��S$�*ǆE���!�������v2�~�>g��أ��X �6�a��Q�u� �dU49�w��MZĦF� 8���i4��+*�"����
��k��h��c��\n�����F0�<�s���K�+�3�t����\��"��B������QG�W��l���'=+�U�+|����X뒹�mFOM�&_�	�����b��f��J�i�K]u����h���M��\f" s¶;�'���I����mW��n}�렾�'KWz��{"t�ɫ��`5�c��Z�Y�H!�.�WTW���?,I��1*G8^����?�� ��o���t�f�%ө{�2{��p��wj��yT�Ɏh��zx���������>�p��igs��j�U�5)���qb��uv�sds$��9<6s��3a-����z��d�{��ㅵ�m���g��� �M~e_)��Mk��v�<"�o*�<�O�2��Bz�1y�u����.� �'鎮t��r�+%<��T�fʓ2S=�ԝ`�B8?��[QBDS�\1OS5E(�$*z`�U��-N�q=�f�/Q��zY�;lf4�Wi+k��\��D9���3AĨ��+�����?��5ظ�mV�jeg�e���jd�$��PB��R�%���n}�+|���=��$�
RT�J�m,��(
o�����'o��sҾ�1z�}
Z����(#��Vu�X�[Cb��V8Z���`��IG�r��S-ۯ�1"o��t��3�7�|8rŦ�=�������2×S2�?l�[�q6��bI����5>�`,��c��(mk��=gF�j�	{C���?FU���U�j�i5S�MВ�u���Ad��j´��g��g�3�~��{"���7 y����Jy;�S�z��L1�C+I�a���@o���5� ����Xxf0�	Q���TK�[%+����G��u|Խ��f��n��a�	Ov
��� µ��O\5�g�h�^$��v�( F�i��ǒ�I籐���+wS9��D~�
��o}EH����r��찇����Ӹz�q?r�x׆�]����A������!���c`����1��F��v���!Kǽ~��c�jC_Wu�l�[.
��"WM��]�3(�"�.�,1���f2$�0]P`w��y}8�� W��&h2p�f��h��{����~P:�q��%6o��Hj;�:��H�<*�0r>�����m�/�h(1g
^;�����]���B��>��8�xC�4[��ʖY[:�"L�:���C]vڷ��j�4���Q�E��eHOH)*��H�TO���/%���j��s���ܵ�IP���x*54|���h��#"�{� 	��V�]���t�G�b<���@	<�&)���M�JI�.�E�ism�"7��k�
�[�Rb���Z���	�� `�Z�>ں8���H���]�d5���f�Qd���#�^u�ͮ����@t>Irp	�ϭ�i v��xP��a��o�<A�p�=��#��z�Qk5���a�X���؜�S��mو\[~���{��S��>	�=3�MF�c��3z�vl�T�:��6�_K��v�Gf�%~�/��4�`jwd_�;�D:\�y	�w�
V~e�[~#v�v��,ү�~©�Ӈ���X�����?-������1q0�E�ZO����=tM������Jj�u稛G�!�J�ޖ@Щ��Ք罙9�'[!1"�!O�X執��;��$�v%��{^׬i��7}���)�|�3?3lJE���|3��ߓ���T6�?Z���t�K��4q^x�2~�JF�'A}���W�}���K������������qf\�U����1zR�C	��Iu�:���:L'��d���àmB����0C�����\�`�%��_�)�3,pvٗ� �A�iqa����邏����@�V�V̭s�}�7����fΟ��'��xfb���ܛ�5ȓL+kR�e!���p�S3�w�=���¾5Y@j��&�g�M��<���d��^;N�9����FH��s&���!�wR�� E��b�x��V�q&���k��D�]%֛.�Rq�V6fd�̑!����P��!�قw�	%#�j���+����z6M\7�Q̹g��${��R�3l�`����U�0F����y����|��Z�6V+��)�
�)�������`�k��}ݻ���9�v��G���2W�$�#��qS��B;W���g�p��D�>������:��rbls��ύr�MEb#���9��xM`�N1$��U����V ��<����<��͵��6��$v�*c����L"�ɓo+��+Y��H�����	�ڜ�pJ[�Dshg+/����I��)��Z��otnmp�Y����L�W����Ix��@��e|��;4H҉!M�`@��@����g����α�?@�"���AS#-|6��pƱf�p~��(�~0�#�s���9hfڻ�ܝ�F�K���:� �rI�v�E�%n����U��u<����(���c`�H��;�dI��R�A��e^�!�S�7+����$�P�እ�k�k�x��ʜ���?@HH�=�H�Ý�nE�~w�l� ���.�>Ҹ�!��!�`�u�:�i���Gwj� ��+���q�E'�k8�J.?�w�E45�_8��j�b)-W�������7�k���1݆ξ��2����Ųu�2��]�Ԛ��P�h[HB���Ei�Q�C�5C~�J�C��jH�L
�H���)��6M��}a�ϒv��x��C�f�������0� ��J�i��%�
�Ms��X��U�-Ny����aB����|�M$��R���x*�蘁)I��ߝT��=翈����,�O���2��I���Qb^��Z'��1�t��2��H�vz����A	���K�U��_Z3&ɖ�6P�˗]9�9{�t͊Z�J���;�kA��5��K]�����d��{p}� �C'��f�7I� n��B/���l0I����oVV�G�2	J����L�Ťk�a�CH�B*�o��X��eOc�<�Vs�:ۆ������ӷh���Ex ��ʜc�C�O�U�w���N��e�T������J�����K����~��f�'����wD�ن��9-nK�:2ԅh]ιm�!�,�DG�k��@e�J���x�f�A�~md����@n?�s��Z��2/D�ˬ��-��|R�" ̷<���#I:1�5�4XYƶD��!�E��9���48�k���	�s��a�����ׄ��>��H��hQ)-!��92�!-�y�6\��L|�]M�1����`������&��!A7Nr��߈�n�z�P�8d�j�,=j�������EՏ��� B���\�d��= �-ۼ 3�����,�Ry���% �bB��FpN��%<���1 �h=� \L>�
M�H|�ɀC�-�#l�����s9I4:����.���i�Wt�U�q��)&]����0�N���}a��2Y��o)Q���z�-�n%%��k���H�=�K��E��H�ͳ�i03��ɤ����� ���M��l1b���S�l�!�Q�=ͽW�R�Z�V	��G������潑�@A6ce�p��<���_�{�3�K�j�"�ٰlgtL3��]@?�c��<���V����O�"���ܧ;��V�>\�B����Й0:��'d1<p9w^�,�v��+��eK�#���t�ZK�B�y��r����	�'_LI.lˡsۢ�z�2y�b_Y�F�?�o0���#���~�3�v�xDb{���������d(�rd�B�i��PU� }3����&ݑU>o 0�MXz Ec�!2�l��--��B `�>V΋�LSM��3��K����P�aK3�=�.����P���r��ɦ�����Y�~���k����f���J<J7ŋ ��WK����.�qZ5E�de�־A[��D�^��FG�0�ҟ���ܯ|��Ԏ�+�7t%���~ܮꑄa�ǯ����]�bN�9��{�O!%J�ӳ\�S�X���Y1�6tt�x~7�3b���V4�J��S$��Nϣz�r��d?uAn],E�k�*s6��e`���í��I����$��������h�Q��TRh"��'�SK��$�$�w��UXH��屏�� �@�X@��&��\Յ�+�P�fjd �,������NH0e*���}f�N�y��]��)��MǫjHh����̩Ph��Z1���,�]h6!+������N�~�ӹ�>5Vևf|@�|Fa.v�e��,��7��O7��rj���7�|��$خ��Hm� �|Ʈ�!��R��"���� �NA
��	j`���"	R�ɼ�ُTn�F(��x��t��8�8��Z>YyIWMȻH�v���7�˓e���
ր�+<���+�r	��K �z��!l��M�1♚�À�m�+�n���������:��dB,.3�X�5�K&9w!�U��ݐ�� �'ڀ��M�=��߹�y��^b���a��\�/�q��:*�Ծ�=�?w�aW	�����[2B�R̥����g�J���&0瀍1tqX�GM�B���ŉX����EG޹A��4Nu�m r>�s��c�s�A�a��gBà���X���ܽ	�Mw1@%Q��^�c!5����X<��f�!5���~�QQ��0f�\[�>9�kAx�Aվ�;���{�|U�6#�����
ʗ���3��y#�����Bn����[�o.im+5�;�����(�
��r��k��h'/ɪk�"�,5/�U�^�~w
�HL<$�� 2>h-��야� g���"��/C���ìO�܋��UO.���V�!��J3u��
��6Tr^2��Xk�����?˟:+/V,�i����wMjQom�Y^�	��ɓxg�i�;<���cC9gz��S�!�)���hq BX�5fF���<yx(>߬@�9�=���B�OHdB6�.κ�M��*��l�H�~#ܠ�CF�(��G.�\��^k\"Ȳ�@w�h�,��Q�ۗ���\9z/%����bɘe��m���z��z�0�a�u�'��}����₸)I^}_��M���֑wo_�ٺ�̲$��d���y��X��=��qʸ���^#��]����PD���Sa�u1�C�ß�8��J�ы#�/��9b}�R�����-�Q���	9n�<y�b�HX�a�^<*����ג͉�%:n3-�şI���M�4���I�4���]��>���@%{,X�92�)"|�ݶVD�GE�L�M��P2mbhҡ����mC2�[������1P:]�>twl��۰�-�}ٕu8�(;�>��L��&!�k掩����r{cTh#����ޛ�x$�5V�@��<��i����؎7m��TF'��"�������r%СΏ!�_q�R(2āx�[^�ūи%��y�d��N�>dpv�UzN�v!��������&��̥���I�C-�'{Ɠ0�h"�x7�h&Q|SCQ�W��53{����ϻ'�ʳ�c|\�bB��|C^���U:K�O����5��&���	QÒ� ���Ա��ˈ}6��д�m�nU8Y�S��ۿ���!@��9\�!tKT;n�/����^"�jS�E \�aV���숫>ls�"�YUԸ˵�ՠt��}��.;�^��5��}�	{F ��pZ�!�y�BD�D��3b!�!��av���09Y�~����K���X� �E>����T"�������Gp��,q<�Fx���(���BEv�NA�����]���%K����D� k�_�o��7���a���2�Gt�e����;`�wKÕ���_Ԁ����h�"$�P�FC���iۃ)%�;?�̃;0���C1���+f�A4��/q���Z��_�ҙ�6�wI��Vփ z�<�������f�T��<i1��P}��-�_��|��r��մ� �")�^!�j/��H���)�uu|�=�,	�7RC=~������)W�>1O�Ҳ�%	%�*�t��"j|u��4����+�V�Y�C/�����NX׳s�'�<t	ebOױ�� ���k��)�i"Y��`����	oqO����<�3�`D��o��ס��,�fs�l=���*}F����p��r�"�,$��u��ۂ�;ˆB����k�V��kRu\؜��������Gr��{S0��lx-��S��iXY�3����PռZ�9)�)2�V׈����W8j����t2c��h}�P�< �;��JI*^>{�݄�*r�qZ�Ț�2��A�ˑ6�ȦR��Xd�T!�%����b�n� �q��ڨ\�)����˻���/��@6���8�����*3���f��^���[|�>�q��iSw���BTԋ��Dnи��5(
8�*wL:\���9��)��i�}����Q`:�o"�жa�EQ�c�ꂱ{[��-��]�]�����#E��^Qiگ�/^��'����n�v�����Ň!FD�6��I�LK)� �~�G-g�\�,�Qv�$<n�Q���fyx�c�5���C�'n��|LȌ�Ʃ�y���\����"B�����uj�'G�^�/wW�(j�yW+mB������k�)��dYk`��֕Unh,g��'#F�̬�� UZN���I2����#�M�&���Y!�|[�Ҽ�¥cj��{��V�3=6d�G�J�P:E���	�{3��5)�)"�*�V,�Fr���᚞�5�5����YR��et�����C-�ߐ����- %5i/l(��ޤ�Ͼy��ո@+rUL0)BI���б9�ڰ�_n��lX��g���L���"E�&�ǮM�ɢ�#U}`��
4%��y�{\û�t��	Ƞ˄���>��`��v%Z�	�7�Z���-eh(�8HG���;����_=&u��b÷�u�I�r����y���&��Mq:Hܝ�`cp�w6V~��=)�����.8s�5�a;��h�"��Z]���A�|�b��%A�?�U{��ZDC�ϰ��c:rX�M��)^�BF�T
ѳ��ȋ�E%��z���xIr܍#X�>#�����k���q=�6����	z2�%��=K�ʛ��X�Hd��̀�� �
�!QʝpvB �n�Ä�E��^���,Q�-Ub��I�$������2��a�k��}e�&n
�!�Y "��j=7/���B��m��S��nv�������_0W�J�p)�29��|uh.��a�d���@I�^�^�3�y[~�q�h�S		��{k'f7��zK�6��~���q��xF��F?&��W����׸��&��&o���lg��	0t�����M�%IoU�bqX���������oȾ��SIS�U"���n���O�'��.��y���'��f<ss؄r���M\%�K�̫����M���i�A�Z�(j��q�h��FO����Tį��۬�s{s�J������}�+���K[�]6�-]b���<����S�{�lrDג�=ud儵Vk�"������Ǟ��P���BÎS�
�4��::E�����l�2����=LP۰/Ƅ���$Qh�	� �P�M5]TA#�{%��������8-��> 7��L�ԫ�*g����צJǩe&������V/qXJw�
��w�k������SMp`^l>3ֺZ�>;ԛ���2�'�C�C��X����ė)!Q[��s�tF�р�54���sj۽��+�<H�W��_Oa�{?�b���!�٧�/�P��ȒQ�:�%L�ᄷYnf����1u=x)HJos1�<�_G�����P��b�2��.�ů�����u�G�U	mpp�V�v�{��bJ��D:�����M���e���͓!.�M7=+��F�����j��>w��qF3m����S]<��k��i�g��	�o�EYׇ�K7�ImO1�Q�����22�ۛX�(C:�Ce6r�� ���C�Nڲ�~��I����N�h�te��٦+�ҕe�څf���YR�l|�3��*<j<��$>Rri�4)l�{5��w����n���~�a8��J{��-+�5F Yh�S��q`���o%�#��6�1����32�vBs�l�^��� R�U�zD��iA�ES�/Ͷ2�!����jJ7;��R)I�t�!�l��P��Pkƨ�K%����3Z�E �+c��ň"�2��ɦJ�8u.�=�o�L����e1�Aȥ��R�Z�C5�^���5:I�#Rq�D�:4t�(VW�a�T2J��i��'1bC�ԩ�7x�N�M���,�NSFn���w4
��^��#��81�!ܵ{�KE��,n�i�R��aY�O�ȱTg��>�c�L�g�HP��n_M*�b�Z�$��'4g�E��x(��н1[4���s��B�Ð����=z=1z� ����	�����������6ǻ��h���ҁL�i^R��1&�ސ|�*k�lt
/i���,g��nNO|H�H��Ag(P/fFG$�%
����E'��� r��0k��_:��T���Q��h�$�=݁�)Y�D�T솷��ba0��`�N����xy�^���q�A���US+��G��DT�wr3��C���<B%E�@��l����;�ȑW�����k���bΨ�P����,��]\S}�04ls�7}P,o�e��$A��`D�8�'�\�>>STy$I�G�M����}���ʬd���%�%������ڟ��8Q0�bȿ�ɾ1�x�<�Z�J�U�@mp�MÛIO�gw�����l��$�h
���C�DR�a��o'�1X@���{�aH�h}�.��'���G���W!�`c�Fu����s�V�ͽ�Cm�C�d  4@�'�5�brK����Lti�~+�f��2J�.�gNz͓+�,i��\�9{D@�GjF�k��ٴ�(�x��;�ݐ?�.�"Y�r�-O���7&��Ä9~��>P����s-���{�k>�� 9�2��=�9��\�~:�TF�D�3����Y9u[�vR����x��F����9�,�}_�ym^4�û���g���1IW%�����]p��d����ؘBz���:�&��dE1m䰥C��^�pbwNڒ���.�n�(�2�y�`{d�~ؠ
ڞ��@+G"��u��C��{����3Q��8֐����dwl/Y�0�\U�̠��*�hvq����H���7��ZZ�T9.��d�l�`OL24`m�o��DՐ.B��;�_z�=��#+�-k]��1�HrWN���c�KL(��m�+�R<�K�$��T{�hs'�0��(�:p�I�s���M�o�juԋ�1S�ƙ�������c|��^�#�d7��%X�	$|���L7���Cy���?;Q�^�;�ş_�����+[���9=�f�~J��.Z�.�څJF�#����ƒ���)�S��5f 5�x`�`�t�q�s2^M�U=711�"�P��@��s�r(	!��SP�OE��81�r��*���<E���r���o<�L�������X�&�J2��0I��D|I�R�P���J$o�6V���7|k:�H:0� <j@?�w�X�Ϣ��{F�(a��u��J����v�pӠݚ��$Sjv}c-F�9�	_\�C�2�`J�B��P��qiD�Nk�0ɮ�prڷAU�@��*��.�b����0���]���ʟ�qt3a���&J�`Ze�+v��3���Zx�	@��X�:�4������#a��?�I�#N�y�&�9JK���4�����>��ҹ��Nb�1����U��֡����E�����e��4U�#hK�3t�������@R��Q��X y��w�3)�c ���aji�����w�7�.
|�w�#yW���Bs�Lf�^�<>hق��$��-�m�R@|Xe	NU��,CWю@�/�S�u��n�F���o����B��z����J�j�3��������<�93�].�!�j�ܾD�@�M�n�C���}T.�tx4�Vf'�|B ��h<�He,-��m��]��?\v�RP�������G�!������@����x�b�2��Ϯ����~?�V�p�T�J�� �	3)V�9
� \꿔���3���O `.��.ֵH��&���&�5^0��]%Ҕk2׋|Nw���4��Uvu��$\��8bT�W	�Ϩ�,"�K��	�%K���_�,��v�x������8h��H����n�_χ�������:��e�}��������q��B�����y*���ְ����\��L~�n$�^�h�Y{�O�Q\�M��R��s������mE.�rLE�Ҩ��" +��Jm���7J�o���X�U���3��=cY�����Б��ܑFe��&��}�y;nSĤ]�)��I����Xʄ�C���G�����ŋ`N���m\�ft��.ke�	O%�,�����L醭��'��iZ����7]�D��1�0t@d��l*W�oa�0�l2t��Q���D*dB*["�<&��v��RP[��	�\����`0�O�p4.�	�W��9@��@�ׁ��{��ě��>�����zҁ��)�`s���W�"�U��b���v�D6�h9�P6��������f5;�d�)Ε	���@�S�v������)2ҥf̔�_����6t���fa z�
!69Z7u�)���!�٦��h�l]i-6��fe�AØYE��1�}!˨)\݅���¿�s_=����l�AR"������bp� ��JR5�W7�-���|���FZ�u6�9��Qg�Y�Z�@z�+<��]T�Q�sh�c��{���C"!��鱎n�%e��j���B%�{q�"5�!XEբ_Y	쩐mU�_��4S�T(H��v�x��'��Ԋ��4j;���Rg�������)��볦5#uai_��q20���VpK�;�|D��;B<�����H���f�>�M`u1]��0���P�.T�����������ş�b��-��v�!N9�g�M�.O��8�t�-���u��q�\b@F�c�[���ꉵ�r5�VT��1����F�%�& �gY�����xğe~i<�G6��.7�T"��Ne�j����),��lE��݂��/��J�������}ꯁ�<��a�&���+k8~"շ(T��dhC��VY]=�e��=(�EB�(�O��|b����2�7+BS�� 9$��Yƚ%�}v i�������O�s���½���i:հ����7��lQ!��f�*@U��oɊ��~��WV�F��%�8Cؘ��2�G�^���vL���G��cs���խl���d����R�nѺ� �ֳX����tGR�zg��G�r)��q�%���D�����\u� �Q��2�`�j��B�&7���H�,�M,A=�tu�+����uF�����yn%s3��!ʔ�f�nf� �ҷ�|Y�_+H:��ٙ\�f�XpH�a|�wm�ϑ"�V")�_7�����6��g��po(W�	uļ�)fޗ�<���<1��Vh��Jd�.	.!>z�@�z��	욯C�,]�&�%�%�r��+������G'ppK���9�C�g�?fS�s��"-��i~�Ƥ��\��
�8���v����F�
��8��ml*�g�t�F��4�� c�^��H����Ǹ��yΠ���0�)��v�&t˹9(�J۰!�q8�Ue�������������CN��+����h��^o�
�$4x2�ͤÓ�N7��8�
���bWR�1�H^���r��v������x�˘ؓuy�\����s�K�ST4V`����En �[N�3xO�^���};B�.�C��d ��uK�
h���.:�\+��x��aй I�� j��'9��`�� }^�[7|��.��^E���ݠ��&�a��B���Ff�-��V脮હ���p��B�F�xڀ�M�<�X�n�E�0�����UHk�΀Wj}�\�yȹeӁ��Ѧ�J�67$	A�_f{�aX�w�\jhW��$���BXgC4���`�T}�LV���Ҁ��AY�j�/��, a��:H���-�Tm�����yY��1hX�o�S�ٻξ�?M4n0i3�<��݊g�Lt�g �>��P��IMd�h���EJ�I��ȾU�k7nt���jbqK�K���J�3b����+��oG,�6UKAX�����?Ώ/l�b�'�*2�K�z��(a9(y!�Ȭ����������m�Bk���`�kJ�N.Z�$c�|�9_ު
��mX��d�0q�n[�ń�M��� @�c��5K���x�X�
�R+IW��G7��[ܦ�K��rD+1|L���B���ۗ�7�D����h��T��l�� AVƠr��\+;�"?1Ų�'>��:�C�M��k!�\;8�¤Y*���e9�(�]M�Ά�xi�a�|�G���ٱ\�#YF�CaBұiҥGQ�؁���8(�'zE�O?]1�}'P�X�G�0Pr��|�D�9�����	*7�����s5�eD�ax�9�g�N��{�km��4��I|M�翗�9�@!$2��/)	�wX-�#ޠs�4�9bn�#mR�"�Sp.��4odK��m�w��P5$ַ� ���t�a�.u�:��1�+Y��{��@����q������c�M����o<�-Ǥd'<�0o��m]����������B#$p{X��0��N�Q�`u]x���+�����3l?w��|���z#��"a�
���B����ë���?����XJ�Xt�� ^��#�U�n=�zO$|�b�q+��0<6aQ��j�sLSG|�S6��v6�kǻ7<<�2����0y�m�����:�9?�8ݞdq��#���Q��pmQ��=�B�X�D��r!�;wZ9PZy巽�ݎ!3oʹ_T#�����6|(���Th}i>Е[��مU����i��o�Z�~b���>XQ��gvV��"����kc�@0�f�M�2e?/�f���"��+?�A��z��Ao���)e��ە2���QLb�޽0%X��l�"n�1��,��p�[������&G��]�)�?�u�h��+O�K_4�4Y�ø\[����}W+�7�R�.tOP��7��[ ��k2Z��f�	�����e2c�����~0�w���W8F��
:��9��$�i>�E�'��\L�T|�:zO�&�:���^�O!��cl�S�UW�h��Ș���S��J�ܶ�.&.N������eY֒zFzn�g���a��^Y�nQF�Y��ഽ	Ѹ'���`��2xO�d5�rM� Pt(��tB��T�Ys4R��fA���'��^����j�4����/)"x�B��T�0ɍ�I�]0�	�!h$�SqDa�C�uW���㌧��3y-T$�1#�ƘА�v����x�2��?����T`����é�7����%��+�ji	�`��K�~�����+�"	��'����Z�MOJp)0\�I��n{��8v�xӦc�����ݽ"9��0�B$��za�dC!]� ���;��K_�Q��|�L}�����<�(L v;�i�	�>p����_� ��b���f����J���,_�w����̝�gWo���;k�$(<��L׼�[J��?���8��F[��y�I"�7�@*n�}�aJ����.�u���A0w�������`:���kh� N��ꃒ�aIܓ�X5�G���3w�*���x���J�P6��{�م�駰Z�~:��/D�g6�\;`ק��5�.�RT�7�)���/�Z���	Ή�1�9���$ǐR�zoP70
P\@�� Id�i�m�+�;rO5�p�M��ä���u���}�2��Hͥ��������5*)K���ۙ)]���睷�W7;��/��٧�W̠qk�s^�,?����;�v�����	�mz�/).��i}<5�C��m����Q����狩e��I��Ϛ
�z�W��������q�[�6]h̀�����!%� BWH���[�3IbȺ�t��mAsO�ȚP�LM�Fr�JnRo��qgjI��	d=�[�QS?���ђ@��z�W�=6T��>�OQ�����k�_�������KO8�,8a�zWI��z�v���l\ړAgd�Ou�̻7��XH�����Z+A�}��([��#���p�Q�C�"���9�o�G���M]�A 1�H��]�AgV �e9֬ܙ�d�����v�w{U�����ő��}e@��=w�A��
�s�ry����q|	9�q��V�z�@~\�`��Dn*����퓋��\�B��ΓuꖕE���D>�O�*-n;�$���{���	0j���ǜ�'�{=��h�A�	[z�5;YRkcz�C>���}:�K��]m��b�ŏy�1�v Ni�W��*�e[�M��~��=F�RFwU�n����em�"u�x,�s�G���MXWJ�c\�N�a2;]�D��=Z�E�$}�[k���*�$	^w�V�	��1��Ř�\��� \��1`�ض����#��L��c?�1�ز��/�]�,�(^���a�-�j�i+��?z;�����:�'*i}��^�?���1�滕^8��'��L�j�kw���V"�#�t��ȻX��+�Ŗ�^h�������ε��d��̣������Jɕؙ�+��/��.��T�9�v`-{L�H���I`��x��I�JRI�GS( ����F���7�4���F-��env�վ��/F��A0(�#%�T��A�2l�SD���!k�}_��-����zM�qP�r�I^��3��s�q�D��^:��*��ڽ�쪩��9���&!�92![v�hIm�����=���u5���`�t\'ŅS���8!���Wl�0P�#˜0���p��yw�D���O� �\�]�3���z\�lz1f)���/��z<��S$#�<8�P%�3;$*�<�J�Y�̩�-<�	�A����{�	���m�@k�U)k�
�	O#�|��C�ƫ��3�׋5$�K�^��=p�����������*^X$���V��#���+�ʅ,�ˇ��i��7�r�X���U��`lR2�0`
.Z�!{�?>D��	~q%�p������;��t��=y��h�zf�ɱrH���X��O*�!�%��;��(�&���w�(�$|���X�F��o(Nm��3>m���5#�I��Cb�@�:�+�f�Z���b039��Z���> O����-b��S�y�W<e0^F3�"x`P��9����mk���t�B���`%v��쯈AK����V���	M�<��ƻ��$��Ls\wuW�V��E\Ϥ��,�Ɣ�$����m �zS���!�#�g��y�����؄�LF�K-���P�]a�Ke5�)�Jӗi�y�q�	y���b7Mi��G�pt�~w��dvv��*a�cx-[~�6�O��BÓ6��p������o5�)��H��{��fں����i	/��C�NX8?��y4q��dE>Ptc�gu';�eEX���%�������
(nԜ�a'���M��t������"X?Z�@0�p��xp��~�L�v >�����P���o����>�����m����A���C=��A�{�+���"������Z���1d�bS�!j���t�@]������1�9$�bv��r���^�Y�S%-�i��KW~ⴻ�ʊݓ�Z�C��zJ�"����[w$��ŕ?�l�r�P3�w^���yy�p��4��J�f-L.���;��\��9iq�J=������J���fy�[F�à�ɟ�m~�e�QI�1���4w�2����b��g��鵫��|��~� ���`���Q�1�1��B�3f�MrzC���3���
rιAz1��f��<���}�&kZ%往p4pp*�V�t���h�㒄mju��"�+د%e~��������Dp;�QR> �/,��r���]�;�P�� ���tz�+o`f*YA��-�����	��*�W�b��X9��q!�e�o��C����O/��i��ո��d�/�m�ǓѪ�ۮ�0(��1�&���F��ݜO��!M*[�+����Q�}��'������qowq<��N;G�L#'��nDFQ�\��Ój-k(�[�np��o��gBM��2K~����/�#���G��*�/5�y�2�]l��,2�*e�����{��Y�L�B[��)��lޢ�Q`�̍Ê����4�J�XKц��ٙ�n_e7�Q�����j���]���ɥbf�]=��S�	���)GJs����Ek�1i��ഋ�NNΟ ���9�[�uv;�0)#�lugQ�M#��|�*H/����]�谞�ʇ T�y�N:��1�u�۷R̒��e�a9�c&eF�Rs(��ɶn�V�O�3���v��5P�?d�@,��C��z��I@��z��o壜�b	b��g�îS5e�{H ��If,c=��AT�ӿ8�D�k7i"@�xt�	Kۈk)�y�G��<ߩ�����|����y���p�ե�c�S#^�˙� #�P�"	�Eĸ��֔m̱7n00_�	uQ`Ȳtˑ2��U����j]!F6�ZN�Y�X2k.��<��;��tU�?tx~���u������ M��.'��K�<"���
��I_���P3E;���m�e�;2��b�y��j��\W�Q�+F�6���2 �<]����_Rۇo�AE)f�}
�LQ,ec�_����qp����3��b��˯����޴�q"�ݻ��_�X�O�d��1u��3��m�:o���4�_�a��!W��P�Au�����B���+L�nEpS��*�
��R`�t��0d��m�wĔ��.W�;Ǜ4m>'���\Kn -��ϦKtnfU�:SA~�j�f:ͥ�9���"q:wʔ�:c�O8��4�uSaȬ:�^=�F�@�Ap�4����"٤K��E0��v9�����vA��!��+���ê�V�Z���"E����VdL���^m��^��灌�ݢ��9a���E�f��O"�L�Q��Fء�X�j�߽?�ڰZ��x'�0@8�IQ�$����~�����q�ju���KTZ*��U�]�WĔA�z<]M'��[�b�j�))�<���{�y�wUP��6�zb���J��J��0+���%������^��D:J�ABs�4�l�ܣ���3��%4#u�>?�+�h��o�$�@b�Ҕp��%��oC+�F����d������M��L�B�5�͞ŀ�N�-�d��DRu�g��^�^.���bDĽ��`O�[`5X"Ӏ�k�O�z`���u�?^Fl���k��v$3�^�m��R��S���D��ETp�P�>R���&ϥ�Ri6>�m+m�y��U?�|5M�|>R$��l�{���H �@�)���+־X����S��dT��%�J��=���D�?q��4ō��ӕ�[��������!io�b\�YR��#W�j���y���	�Z�(`���{E��#�>�ѵ�{���q\15�}c�Q���)b��_a՝���H�b靑U���l��ǒ�U_��I�{�|��x�/-̖­��OP�� ��^�w���Z���.e1��rI��CHqK�z����3t��Q��TWvV�p�35�j����ۏuF�N٫���U�G�=�{DU�$!����z�k��_u4!�%W켑]D8������[N��`O�Q^,G��yO^�Y�=�)Q�4i,�$�!I�7�BQM��:�V#
�; ��싂ԉ�$E�9&��[X.Ar�vר��{z&�#m��-^�����*���uς�AI��R@��+I���4rHI6L�� �Qf�b"��h�΄��l-_c���͸��N��j3���2��'6"{�/���ˠ�������1H�}�(��_����r%	iH]� ��1�#��(V�i?��wϤ���!}��)˓J�w�z@��[���}'��l=�� �u�C@M!�k��{�z%5?��ϔ,��J�lq]j��.G�� 
��ICn�̸��i�f�	��x7}���~n�Rǟ�p|��r�ҀA��,˿�i��*���ow(�l+8ac\"V���3K~D{6�ܗTm�	��b�A���0a�N�3V��+7|�u�[(׸^������#-��㺙2	��a��Z�G��R3j�Fޚ*t����Ոr1.f
�B��e�Գ���QR�#���b�p�^�����:�1���y��?�/��p��i-� �P��-�ed���+�aNG�G����.����NyJd� 6f6��x��j��6�Lsq���^���8�R��������ȚݙGX�t5R��;<��O��B;�Zɡ��@��E���+��RĎu�n��=�S���K�H :ZL���(�H*������C�!Ȑuwpx]����@�c�e�t,��Ww��C��mm��C7��X� �p�a�C��f���K�U�ӱ3z=	~��-߮̅��T5�s}v�Ek���/p�u��4�^�#큯���5?j�zsp2���jN����}o3����o�T)�H�a�O��#�6O	9�c�l�>W�Z(M��8ƞюg\�KB���v�� e�mq�.e8[�cn��_��|	�:�/N'�Q�Dp�k��A��Y�#�����'����p���,����P�3�|D���o��͔p�K����ՠ���7`�o1EӒY����p9��Y�X�gXR�"�\i�n�; Aݱ��Q���I���R�J�:nU��>@�\X���Ԅ���IRm�s)��<������sL�[!���� ����X�%�[�
ѣeRF2�R�����6��P.4�54+7X�T#.F��%BK�t4�Mי��Ђd.����u������ʺ���?r~�-������wA�#>?�"�*<:�P�9k�,?�j�w�)F�Ț��G���+�E����
�G!����(�=� ���D��Is+���������}j�b�k��5��0�u����ȸ���7�;ݻAP�*/��j���B^@!wƫ�^�{�������Z_Þ���[Ԍ�`�(-KGz�C�A�6[��F"b�TR�u"���� :B���`��:���ف�0�}_iHJrk{G
��<k�,�q[�!��y�_��2)�h����=)�!��j�S< ]R� �W���8T�@ܸ*�p=����6��Z��ҶX	F]��ߠ�d�:�yH���ชr9��~\����p|F�.��'7�֠OBp~N/y�̳��es��K6�����)�n�/GlihÒ\�	����/6u�T���{¨�45/)G�������_�9��mc7F:)wMt2���82�O���ɚ	��c9F/m@��n�;�B�O�v����=�m'�ۈ�H�@Zw���;p��	����	R�`C�8vK��/EJ�g~�̂��f%[�]�B5��GRUΪ��4���J��"I�۱i4��"6�=M�Է�;-�]�&�cۢ�l�$#����%�ν����M&���@зeVz���M+,Q