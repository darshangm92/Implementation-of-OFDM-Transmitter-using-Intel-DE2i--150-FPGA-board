��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����軥�JƆ���,����TL�����cߣH�ϫ�о�Vy��/B�h��I��|�I�%=$Q>ߝo�׬9O��7�ٶWf|�$��E7��x�AO�&BGFYHO\oe��V���ન���*����������8��u���e��fA�2TFn��$�U�p�.�J��?=��Z�PClJ�p�pxhΟ��<�V1�Q���o!z&�"d��m+���ESE�	�<�f}]��q��9np�i7<(��6��t���#E(�F�����n���-U����Y̺ ���Q�}Zm���04Zȭ.|�푲�ݝN��h@P�>���/2<�n. J���O P�6ֺ��X�"�����2�&%P��Ky����h�+pdx�-E�b<p�Y�%��?�i�J���x��r�15�vdX�*�K��(�͹{��h�8��1i�=���G��͵L�5@V2���ls��N/��G��܄�kT�wA�U^�Mu�@s���|A#�V�}_�>Hg�'��DH��SP�N%�U�^��;'�Q���Y��ˉdne*0�}QZ\��3�,{'vl
��8vUrY�z	��>k��)��qO1r�W�T�
(eN�_��1�%�1@���'l D�2�mM�m��X3f��|�q巗x��í�l�]�H����\��n�.�_���^�\&+�9z�]"�_��ZM��@����kW���ȶ�?|��t"��� ����Ɖ�RLk�ח% �����gt�Y8��pA'O��fgaٌ����8HZ�A�S+8m���b���t�r)���W��<�V0͊�-*ޘ�q�n�нB��ѢVH���|/��|�s�sIa1���5h|"Y �f�ީ ��$��g3�g6�������,M�;A��<f��ce8�9��b�̋��6���)��y=4x���M��RfZ&+ӡn��@Zy0=3\1�o�R :��.A�j�K�ܑq��V-6��<�z6D�7*�"��v��i���~�R1:}����4��;e�������웂l 7����Z��o
e��u��W{*�����@���(���͡/�"�v3���T6rC�ikL���Z%����v��s��5��,��Is��4tL3(�=�w�<3\��!��j_�h���������+zz�+)e�]]�@ў�X���Aui�}�����"7R��n;�Ԏ����>��\BJ�l�r[������q�|�9����E��bm�D=B�xB4�K�1'��Qv����Og��T��R�aW���`u~D�ش}�^�8��o%X�\]��C����Yl�e|���B(e{�kx�y���	��s��(�\1��ͪTN�4^�E�3܈��7ZQ�*��z��풙,��Sd`�/m�zY]�a[&s�}N_�6�tn����^q<"l8v�X��"�n~�o�{H���xX�c㠑�y:����;�$H�E��OH�����Qd��_m����9pQ�!��R�����K-^�L�"2��\��,��2'�s������wH�'a"�>�ى����za�F>��e�M�5)�����O� �ٌ��=a�����x��9�0���ĩ`��c؈~^�1k������V�/������}�+���]������ɢ��q�4�V��H�}A7���Ka:_�G�7�&<�= �`�y�b6�4kΎ�`�
�馲��>D)�R0��!�Ќ �G_�?�g��%�uO�a�R��1=;m��Ϋ{��O�uM�[��5 r}�s�E�{������`e�����W�����BN�w,�9���13��fc���6�3�JǐBy��,����D��y�U��\"�������ew�����(�E�_�Ꮑ�P���H�"�:���z	#�(�^�L��lW����M��C�#|�_yh�!��w�D\�,�O����@�B��ɡLJmo˔��ڍe ����C=���9	Ɋ��Յ Fh��U�Lq��I���XcHMCF��m��0��=�h�gY`��+���D��;���zep`���z�#��]���H���1�H������Y �m�؍�|���JI��Y�-�Ux�K���D�T���~�z.:��M���վC_H۽0ݻ�jX����R'Ύd�p+9Ĩ��ȉ� كHw����i��GZr�t���3�Na1����]9g(l�#�	�@�"��5��h����T����K���M>��Yk�_>�1����h���߯��1jc�����������@^�$���/p
i=~���Џ(I#�]h����j��k׎��z#ԯ��5��ΰwLn�|�l�?U��pJ�S/x��vR���|�c�H5��k��DC�@�K�:;ν�"k���,L�H�����p��UOg��ωP4���I*��X���K�{�;��!$cW�	����� 7����� B����fi6�������҃m��:�
��� �/��l���B���V�˭|㢉P\�(���:�������^�.�U㓗·��A��ҽϠ�Uiu9�)L�K�5���7��/L�������u$q�����T��Ӓ!�\)���"� v�01�U��V�Sd��i���u(r����ڙ���^ph�,c��$�F��0�s;&���~e�*Rpk�@�n&�Z@���Kآ��C,���a�D�pq}s!��U�u�S�c7���Q4~݊���1�Q_�CS�̯�/�@��U{9d堲�u�|��Apע�I�3���@�nQ�q�)"U���wY����|�܊y���p��4\�G|Q��η�,6�#�J~�ݝfb: �ӍC��XpO(�}p������]��g��2�cU�d��F��:���D�z]{м*�䵈n�<q620�1���}�����l�ъ[�n��`s\��Dx�����Ķ�N�j�o�z_�����Y�����#Bj�-\]��S���������B�L;�Ѭ���R�Gi:e��GY���i�_�V��Q3�:�iJOe��s>7�ƃ�?��Ek׎��+�Py�$���:��D�Z��Kl��Xg
��9���)u{�[o7�Ͽc*A�����<�e��kr%�p<���F���B����B�Ug����i홂%6��$/���{�������NG,����E(BK��0�9�lg�*��@�Z�F�� 	��Ri��n�]bX�ES6�DZ|�e�=|�1��_)K��&�"�Ӂd�1��3�%dZ��O�$��c�M֨���&q���&���=J����ZDs!C���U�4p\�����\+��P�?�d�O���S�_Q����������8-2��I&��^Jt���3�9�$�v�h\�dĀ6݊��{��Wݖ�`5��%b�~-h4���p?���i���M�?M��&	�E�gT�&O*��+�A��F�͔r��Ku�*�LF������e��̡Fi��N�?��i"��>ō:7��JH�}4(����2� g}*Ė9�e��d��ɹ�w-\g=9�_(���7��U�/��5(�˘�@N�L֟���~>{�,~�_c��OIR���l%?YEԒfI�� �`XFc��KC����/�n�1���e����F)q����F�sb�i_�<�d���m�ދmU��M��%|�J�hhl�[�����ה&���B��I�Hz�.\Q�K��o�RN"����O;r�H���e�e���c�&��L��?M�:L��gQ�_K	�Ʉ\��~�%��S`<G �?��R�4@ߢ�
�vv�$W8�������6����q�O��`{�k'Eh��n�h@�x�}�}R���1Y4[;+=5���W����Q#���� !�������B��2%k���RhX�m����-Z��E�\3�O;Yo�w�-��;\T��ݙ������2ښg��G�r��/��Fi����2�ܟwe�)⺅�]�lu�  �����$7M[��!�8��X�[=�Y�
&]Ϥ-Z�A�ۆ�G�R�u��������23�K4C��S�G�j�i�FuVDz��^j�U���Z����~[��0�%�����5_�vyV^^���2C�{�
Ǹl�TkA%+E[�[c����u�(�i>�;��3j;����??%؁m�'�3i�x H��U�%o���EkF��}�K����qzL����q!��HwF/>�T�JBDT�Ox�d�c���ҁ�3d������I.G��a�����I����B�NΧ��]�e1�HA��(�R��<�Ì+��#"SC��G��#��'j�e�V�}��sɵ4���4'}�Wr`@�a��8Ƅ�VSune����N��}��ŏ���L���c���Z���A�Y��+�ڃd�o:�:�/��u�|+s����Qw��'�8ʗ7w��l���`^/IA�D�ʨ�釓�jP����h��{�,oMw7��0�6"�.����C�R�����Df��Z���}O���g���D��V֎��C%�xȈ���R�պH~�)& �z6P�G�$�V�Tt)E^$R3�V��D[*��9�h���5�,�w@ ��{��*�Ѷ[��Da��ύm<EBm���
���v	qk@T���zs���C��ja� ���&�ؽD'JX�(���kc��
��� yS)اC� �������_����|d��)���m�D��ژmDP���P9.���vio�+J)����Vps�qX�W�����9��X�ᙦڐf���mQ$8��x��Q����:L�-�G3d,��lL�j��#"�]��A6�i��3Uf��>�a��
�2��-z2n��f���%�y*�v��Uy���d�Ŕ�9�$�|1�9vd��E�#i}5�50Y���d>�%�0���Ӊ����Oܑ�5q� ��-���9�|C��l�8�kѿl�={�Qq�^^�e��W@�=<炓��h�4;��Ю'Շ,�_��E�8(;I��Y<y�o��U�7�]
,Źy�)qA& �Wk9�/7�Z�δx�����'D�P6�9c+!,f$���'��)�@~��u$�v	�����1�&�߸UZ4�W�����T�E�����9ۭW&�a�D����A��)E3qoſ�+?����X4H�9�?e|�D���Ϙ�#8����w�"F.�|�Z]~���=3���7��t-50q��%mmZVܢU����~}��\�bA9S����2��,��g�Z��M���xP�0� �Z,��z{+�:�$��:��Hf�A����+.�/�H�CG'FB4�B�:��}!�Y|v�# ��,�u~eL�ĉ�ͩN�v�7�������(�P��;�j>O�2<s�)`�����ZX�����3יע��Jֶ�qЏ]+�/updK+�G�`�o?��^�O(��Bnf=���2��v�Vg�λ�y��ƿ�-���$��-��~�u	B�,�̇�@�Bz
�wd�5����y��w��)d�J�v�1赇�9c�P���ҋ�&=fBkJ�K�(�� V�;�-�Ha�FU���gl���P�y�3q0x����n�,M\�ʎ����Έ *��<��p�j_���f@wB�3~#u�D����?k�c�k|6��EG`ʩ�ʜ]%'���g40<t�緋~�b���]2�\lOK��r͵	���g����t�*�͈�Y>��Y�\ˀ;x�ݾ�U+���7��*���MC�Ĳ-v���E�g�\��	���e�~׏���6�
�J5d���BtH;�\Cl5R��6r��΂.lr+h����g�L˽H���bD��B��K���&
)<^�%�Js��*0���D��3���9n�/��i;��'G�[�dw�,�膂c/T}[�w�T�I����h�B���:ɍ;3>-_�.P�i�s0�͋+Φ��57f�&
7?�38/R�?wR�bo��c�D�he��c�v���%v��&�і�Bv+�/nk&�BC<#h!�ѝR�n��C�S�)�8��aЉ�D�B#���9�̾k΋�w��PJ7�4�Y;���d�m30�6}=D��2�W@������Ε}A����rԢ�o��ҪW�����}b�R��-�hLN	