��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����ﾍ ~��ąo��L�N`�	?|�,�r��iYHڞ�T�/�[���uİT��j�	Q߿��pa��zxX�Ӥ�T��H_ދ&-\�V
���l$U{wص����F�>ܼǯ�HW~"~f5U����s[���~í-�P]uǘ�0�x�,W���$uDL����e����[D)}*z�����Ȩ��~0�roA��:�F7�g]Id:����_�!�rsKԝ�*m���S��(�
�'7�Qe.�w�"W괼���.QE���P��e�E���Eù��Y�)��X^�2���j%��U���V�X^�ig��el�ԗQ1@��Lv��0�T����$�鎥�}�u��V1�����ʿ���@����9F����2l��%j�&/���]fO�{̵�u�#����#�{�]?�JV��6�TE�ɷm.�`:Ʀ�M72p��1��IW�J�a���{C�#�隳#�ꍭ,R�� �.�zl�ܾ�au`�w����8f�̏U1[i�T��li	�Nh1Yؿ6�����s�9à&]y4t�����%��vDf�$�3kZW�=D��:�f����������i܊��5+���ng�б%�'Y�"J���K��~pc�U�ɦ+�3b<���zRˆ�3����eHn�#C���4��h�t�,MG�6-���B#�6=`!���g07T��X;��E������T���F��}D%<��"���I�5ڱ�uF�b�\�p��]?I���"¾�oڬ��m�`�2�)	;�� ��l�v_=��*��FFA��`!������"dQr̀̀��)Y�\^���UfʧI�����lw��X�!��dЯi�r�"��,�a�I������&%!����.�I�Rb�b[����L�2s�Qڲg�9k��F�c�"���oBFt61����76i���At���2��iN��-K�`+�T���fρ�Kyl1�\�W��MtrS�M��~ܠ�tg�ZTJ)�ߏ�4���Z���k��G���'��ṍ��v���%�P�b��aI���*v�[��qhp��&�����H��2��`GF���)Q�!�5C�!�+*�-[���t��Z�*S���;��A=C!7���䄑��@�؞��1����Q#�ϻz��jw�
Ц�s��~��ަ�/*Uʼ�ɑ=!��_�� e5j�2;8��0�U�u@�:���[���Q����Ī���jm�+K6�/XC�hC�ՎW�\'�!�J���y���p/"*�r�� S��Y�(�Un�?br�
p�n*�=z�(��T�5
�}W�7�Z��@GG��b�Y��5R���ԟ�i����ݣ3���CqTh0-}Y��JC�y���Y�vp��r�QGӣp\Q�V�_�G�`SW���56͂�j �B?7��6YG�U��^�	!�8�Vd-�=/@Ϻ�=�e�0�. ƞ�EX�3���S���󣷌\���$e��D�Sy�e��b�.0-R�F:�ڱѠ�� �˥���뵌%�G�"�?6ȏ�l&k@�=����Cw�c�29�.��9+#p�!�I�����^��i�a�7� ;��/(��7���IZ$��)�_�R��lԝK=�P����H�L�D�1��Ց�*��X���+��s�q�*o�����:#ug�33�J/z͟�U��>��PYt�Ϭ ��ZYD��<AffN�ɩ�m��-\.�>@��m�Ts��^���T43@U�(�����'`��h��V�iX��rLN`ʈr�A��h�[�
v֢�>���b������h�F�hf���f��"�E��G�����=�<+��7W��]��R�e=T���E�Kx�
o*W@OFcNg~RUٍ��s͸5p�R[�EF7giѧ�_�Z킉�sO���bpW��@x�������Z���ByIs�6A�t�(D�;jx�
r�������=I. Eq}�NZ"5/�E�kD~���$ �K��(}�6d=�c� ��Sԑ.�^Π��� "ġ,.� S5��a:kF��� �\�޺X[����l�ܝ�dY�SqL]�G�㩋�1a��P	!����c����"$�}����V{�7ֹ@R�Sᾢ��-���˚񿚸���4B�Tk7n{�di��:�Jh�F��{K@�$��z�-�/���hTH�XUYuվ@��¡kh[r$�ݽ�1�@����m��C����.�����$w�9]��n�)%S��z�w_C�k�g�.���3�������R����Ps��Ȩ��u�۬�J=4x��"�C�a�K�^�om�`z��)�׷w;X�@��k��,[�A�'�)��W���ˊ�7�b�|����ڬ�mK�a^�ʶ��-ae��T?TMhK���-��ŕ꾹��a<~!"�w�g6��&?���J��%�����_�������x\d�i!O�r!O~��{m���U��Ďۇ����T0�U�cَ�99KCa"+{���?4�H�T��\K�Jͳ�;��o-E�Nh:���'�\����s"��=杩G!{��l,�\�Q�˫&��;X�j����N)��?j��|�����F-?H�íxm��٦5A��C*'AI��/�D��y�Ij#յD������hb%�s��I�&
6�6���yˋ���z�T\���˰�<�.�-���g2�e��M��k�b��SvT�/n��Tm��L;�|=`�)*\��B��"�}"�޾�/�ޒ�����j����'B@��9��#�T|*C��%�N-X�K��f̧:�����\p��u@���7E-) Pp4#/3�M�!�H���d{��4d U@C��ݰ����L�uے���|9.6��W��ܴVq\���T2��5���3�g�<�(�=ϼ٨��i�����jɩ��N�h�jS.(���� �ei���#�Nn�E����Q����ּe��ޕW�<ƾZo6W(I�=ۻ�BAO��Y�Mv�[�_�����!pc��Ұ��B
;J���I==�0���T���bc��1b||�۽!]5{�������Й�r�I�gi-����TaE)��O�xl���D���E_%D��Tp�[������f|i�=��	�T��]����o���忠��&��]���ū	�T���sB�d��� h%N;��*�ĳ�z���r��/�p���tr����������U�ML��3����x,��Y^op+`0�/��ă���W"��[k�Ƕ�r���U|��z������#�:�I�z\��reN��d��׫�������H�K)������Q��
��=����4qa�g�6�d��#��t����ș�p����'���;����F�oh��û�2��j�pZ�&��k�]0�c��ou7gj_3����|""�X=H�?��2��9�(���Rͥ���,�] Y��L���x��=�PoW����]��`b�^'D<H�ZP`���d��g�حE��o��Q�-�f-�7���2�ƺ�s5�&�d�^�yk�5R��:�1��	�ҁ+u�#�j;���}��0�`r��^�ǁ��$���O��d���yGB�P	>�!��?_<6����-#�3eB=��r UU��΁�~���$	��|1j����*T �fu���r9����e��w�P�_�5���mZۅ�qS�L\g�#���V(�~a��mkT���?>-1)�]h��%�y��ӡ#p�&V�&�Ԓs�KJbX�_�p�q�Z�6����E�]�N����d�ލ����D��5�JA��3��e�H`�RW�����LB9�Un<�o��q��R>O��V�U�Q�P�*Ϊ�3(�ܾ8�}4H*ى��i���ǽ��h����	-��r�=Ql=����`����|��R�Ԓ���S�/��7���H���x���6�o=f��qŐ��_�7YQJ�juz,$�8*��_`X{�{(Z<�j���c��M��)���{�r��2��� �ϰ���ճ�7����#x���s�f k<W1�XL�	x�Ϝ��V۞����tc&��8/��_����^��| �������pu�w�B�������;t��Ao��?��Uw^$�� ���>�AH�o ��;A���/=���� k߀Wد�Cq��Ś.I�\��,�X�ile�%��N|@�� A��.�`��nH�W�@��!���VPN_� ˑ��q#����h��l��%��"]�n8��IT[�^�\Emn��xc1�ri���`��i"뎟��SɡA�2�J]3��MO��lr���G2�"�s�?�(���c�'�V�E˶0�\u�\fU|����j$yi�g�6!����U�X�Xp���K��{F�.��X�w�G��Z�l�ä9��v,[���Hgod�M�Rje�
���,	s(E�S+�4Gч5���gf�h\����U�gS�@��VL~l�2!G(�6�8��n�2����]��1g�#�LЯ��RM��׍�}2e�1^�P�
h|H$cb���X����|����?Vr�4c�.>wFY�e�� P�qxb�J:
���h��5c��D����[�����2�2�O���G�uh��-���;BῈ�~��<[rp�K���6�_3�fB����ت��Y�s:�R�b2{�\i�	�*�:��~��Ә(���?H7_��ޱR�X_Zq�:�ϚM��n�����ࡧ������o�t̕8�HT�f�P��-xit��خ�`����-���|	d�����k0Ǉ	8�����ܩ�2����;�m&Q!�3`Fj����-4�7AT����f��~tQ�ȭǙᬋ�q���p� b���}R����!1��ne=��H�LS�%[ߝ3�\��#�����	󝙋�g=�����w�ɝ<nh�q6%rD���V�ML���i�+쨤�����2#Ԥt���_�V�nUO�|��`�'J�ug1�M�qs ��$��cfwcV9z{_�"z��d�N�2��#�t�x�,ϋEJ衆Ur��&�IN�P���莄�_�SZ��:�3@��nFe�d�GH�.�����[,g�h�{)~���"�6�}�Ď�G4�Ul�`����t��j�������Y��MP��Q�o3�&T��)�Q�B,9���{G�%�l]��ܿ�I�L�����7u�"��jD�~�8h���La�u���O8�<�ơ��Ĥ��!&Q�+���@[܎��'>1�Y`wy�BV̂*�DY�cy�@՟�@�[m"�A��@l�u�H�>�������-�F�����͢@����k��棜�ὛW~3r��(�H�bę����F� �������̐kT�=�qDPŞԊؔM3�h�h$���Eb�����������6��Ɓ�U!��>�3IW��p7�fbcw��܉d�"�b�O���U�"Rj�6Wo��a0��l\�oóo��E]�՜��!�T͖RV�bSzwb4�9�
E`�س6Q����L��Pm�F+�e��;��0P�C���P���3�Ǡ��h��=�'��������@����o�o����Y��u]�D�p��)��-N7��=H�X�
�*5(���W�TnqT�p���	�c��6�%�DF���u��T9�0J��۩��H�6��w���8�ؙ"{��I�#�=ߖ��szϞS�{ &��du]�?2߲u��M{��,E��DKK6X�bYFׯ���2WW�j��l-f�"�
�����VH����9� ����~��H�w��0�&�&�֭!	����]�0�븵�#�[b��h��2�,��V&G���T�W,��w��+��&l�s@Bן�%�YT�Ki�0�eft��o *�O��^�42^��}��$~�
�G{4��(Ա]�]��7���5�_{V.j�5ɂpz�}w/��Ӂ�s�� ��d�c�����1/]b-�ů�y:ч񑩔��RGb�FL�5���<a�~V��A��>��8�	a��N�8�b��WD�Xd���c6�GZ��AP�H�Jղ� 0�{.��	������K�煙�L�!H� ����d�5׉u�CŤ�� �C�U��h"��ǋ�Ӛ'̄��{��ǣ���B���W�B���F5�Rk�)��
/����GLS��fc�ޥ���:��Xz�i$�������\5�O̰I߇)����A��c��?p *����IA�4ZL��.�#�n���� �,Ц^<��Гǳ�h!뙾Y���'?��$�R%r��B��GQ:�L�ؼ��?�>���\��W>iv�N�g�1�k�נ1i� �ed���o�� ��/z�C,�u��܀�@5vD�}����&�'�p����U�ne/4�h6�>7���5��^����-kvɎ>�] �f`��,^ȡћ�z1#؍�Mb��)��fC��YڨR���J_#���e�(�����v[�Q�V����S���aۥ\c���Q��lw�m��OPuEc�F�c�.Jfm�Ii��b@.�p�y���3B3!�y+e�����$�n^�ď����;�^A����I����a�ϷN���4j��f�-��ޞ��;�m��7!M͕2)
�'��y���x��|d�"���`Nܛ�X��tҴ+�ʦ�tV%q=�R~�X��.4 �a����7 q�8hC�h�����v�	k/��`��Y� �Lӎփ�7R���7������x-LՌr��=l�� �j���	c4�p�\	9Y�&7har�C�ڱZ��P<��Z�FҧK���F9�сߞk9�I��zbN��Ġg?�U~�'�����B-:���G��"�k?�G�	�B㗫K�Lȏ!��E���s��p	c��W��/".$�XɎ���\5����a̟0����Lf�T�:�Ĕ��aݘ��
��XT�Wɣ�tKH���F�_Js;�x|Gb���`�s��&��<��+s�A��G�b`j��nq���+�y-�����I�S'��tq��K2�X�N=d�Q�q�9e.���e�F�F�}�L��0�;�XF���"�y8��n�M7>Q7S�t;:�����(+A@U^L�H�2��=�I}k�h�$8c�p�?�_�/��ߓ�#�K�T:[��E��*�HBvW]��p��- �I8v׽=��yG艶����t]ְ�6Gtuء�����Nr��Lb[ޤ�l���3�������(xB�u ���!���Z��a����pP��|�D���oP�%b˗�A��}����?:�Zҧapnш��ǊV�ؕ�9�� r����j8w��+;S��ٚ܊�)����U�]�y(^����A6�����%M8~�r_hP)�E���?��1�<���"M携\cM�&hi�����I���+=NBm_����`�˓hM��d�4�[�
�cmq�U��!N�IA��[��J�!�zJ곆B�s[2Tv1&c��;6���;�[�gq o�*!hy���Z�3�7m�����[����V1���E^v	O��uH�A���\oZAn���9Ii�@����ԛwen��2��9\D4	���]?8 ��m�L�u�x���V�����٬�ɩ�&.Z�"�\}V�ݟ?n�D6x��9��Ta�;�����d���Y:�%:ȳ<���.��z��[?ab
��b�2�Cz�<�!��'��N���d���M�HE�K����LQ�	Tk�GX7�5��Ng�YW�"�Ô���P\���z���5���t���?F��G�ʈ� ��Ô��i�rR)T�c��X��K���%�%W�t��ϯ@I�F�>罫u^0ήe���*E�=ٖDs_+�f�Y��{Ɗ3ߋ3�uP�-��)�ˍ.# �:�b�����V�M8}�6�?Hz�XI�*��^fހ��
�魡�Y��U�,��Lե��9%廬-dv�|���(8���w�Oӂ�э�'f$��ݏ�k�d�����ܙ�"�h8(�lJ�$�j�Or��tfp�^�a�PQ���@�(���k��vv�*�*)nT.˼�3�R�g���\%��>�ީ��d�n���yF��:ݡ��@���PN��L�r��7v���/9\���p�*��	d�C_O��sˣ�U���5�����{U�O�b����E�P�O5�t�WlA��&��$]�7_T�3�O��.�|�Fc���r`���f%����rp3V�_c����$N���g)�b��S��>���.M@\���!��X�b�4=9����a�)%ȣ�ޘ%[9�yMn��k�%ӣ��JݞY^�.r1�"_	�+��//����i���c5b�A��Cŋ`)%�^X�8P���y�ɨ�����_ ��?l�s���Wu��JG��q�gY\��P�j�:���c���Ꮟ�ݴ.�#����I��d���X�ZWܨi��`���8k����Q�A��XŚX���-#��=e1η�CV���	P���O�����Z�DjACs"I�-�9V��gw��4MQxE4�{��)7b���́,�V�u�8zyg�Ѹ�`���n��;��y}����)���!6���r569����Ps���� g@N��76q�% "�V�w�,���CX��q�F[	�e��!�/&��Z6{^�o���DS��{91uw��c�D����#�t����5[)Ge�S���,	�~���#䜪wW-�v��e0��I+D�����t�CҍBV���~�W�^H߮6�_5M�.֌�і u��FO�x�G:X�/�A@��&��Mq�7�sA�ψ�$�;�གw��wC�ch�Ԩ<-���cI��M��2�#�&ȸ����V~�/�����C��_�,8h��t��m8FD1��]�m��[-R}Q��J;?�eF`(nbl��;���@z%JZ�FX��$�k�)�l�Ja� �0E��x�M��s�溬��S��&�v� Rv�'R�r�����Fc=�y_#t#�P��h-�߲~g�S�*4�����%<{צ[�"�E��boEP�b�ׅ��ińҷC�Q��*�,|���͟zVR���)��e8��X!�<���N���b�U��J�����TPd��l���)?ͯD�u��V Zt-��+���Q���`b��%���{h��!�ِZ;��W��78����/�?+a��/=jxT��;�D8嗃2�R��6XS.x����� Ua�pO���P�_�^�y�z V�>������������˦/�^T�	�Qk����K�?.]_�]�t>�O_��#q;r�jbQLh�_j{��	 DK	kt�B~/��j��ob�3/��>��Ł�=f�]/{�,�hD���� �[�q�Q2 q����ɕ���|�tS�mЬ�QM��?g	��*��Z�h|&�D��ܵ!�X�T�oj��ͪ�O�ԭ�����^��E�>��Ԟ3�������҄x�D�[��f��4?&�6Ȱ3X�B�l��LIfc}��*�G��k�=����M�fk����;��g)9�������Neh@�"�����I;,�tS�2��]�^�]ƌxF�8{<��[�d���Sڛs=�,�h ���3�m��"�u���O�O����1�:��"CD?��ߏ��F@l֌�qo�H���w��z&T�ޤ�h��d�a��&����4A�!�r�X'������NL� pY�}��h���h�)��]�ZM��R�>����f,W�GN[�+���<��1n��(	��nk����x�)��]�O�<�[M+��$l=RJ�-{b���z�v{Wc��b:$<eA�E�N �xE��F��*M?}Z�I������~ChD�M}��S���j�s'������W�փ���*��d(�z�@E��N I���X��[��̒�e�\^�k��vȴr���ރ@��
&���2ˁ�����Y���X��-'���Z^�pca���i7�,�$��:�5qJp�m���_:��e'�1V;���&�c���7���o�$#,fgH�p�7)/֓���o�E�O��JU�"�	�v�G��ɞ����/V �M��
�d�i��5��G�c\�k �֖�r7,'#��I�:&��!��"�A#c&&~�T��>l�0�����ݽ�j�������U�8~�k�>��'�LK=1��\���w������m$�q^���VI8S�Ta�. X؎�l�>[�p�ߵk�/��p����Zw��:;N��K��4w���<J�UeLjO�1�}`	o��aR@Їdm�nZ��
��̿�ҜQ$�K�Y!��Ok?�Asu���l��U��w��ώ۸�g[��[�]���t��ץ��vq�h�HG{�Ȉ$���a3��Ow�="2����w�4�5u'9���Ѯi�eK-�h>]΄�t
T�g�:��r(�Xl���o-R�b�4���0x����B ��~���C;�=��!HǍ�wn6�d=�SёDM��O�`�\�����AWZ�6ib-�{���k��p2+R�a �^���]Z�r����,Ы��A�8yL��b�A�������|�q���j��Q�/�o�- �A�8(�Ӧ�ƀW}�c2��:B����S'��a�Eh��m�*�����S���A�����pj:ɷ>qc��h�[I�L�⛠��.�x�]�.{ê.���(��E�)pcm�:Z~v�d������=&BD�>�����B��Fy��\���" ����AG?k�:'E/���<o�8z�)�C�L���=R��=b����eB=m��Q���0_�i+]ԅ����(k�E��2���(�bNi�{�g�_�� �SLC��߼'�ʫ�KHy�nIɚ���hY��A}�^���)a�|�基]�v26�GE����8{�ۧ��)�,��^�QM�D;����׋ɰ�����۶=ޛYc�����p��2v+.e��f8�rd6b���@s !�O��F����{�[][u��Mǧj'��T�@�mb��޺6�8Kv���)3W(���c'�'4Qq�^��z*3�X����\U� �lr��oq��9�鵜E	W�:�T��'I�����;'��[���#D�gO���m~���|(eH�W+
ҿ�H�~�O�a��I_ ��	��?-����r���;�,����`�(WT�k��u�č�Be��_��]�	p��PC�6񐿚x�Q-������� �wGf�pV��J�W�6��W�yr�H���U�u��S4�i.}�CU.0�Q�{�TD��y'C��)�� �����p@��#(�֌���z+�*��a���Y��-"�x�ٲQ��!��ŘDᄍ_��y�<�&�H�2r�2t
x�w�@C(nB��_���5>q��KA:�qM��R���\l�$�J�"^#�#�c7�v��~��������,L�F�r�G�\�l���E�@8�>�I�ƌ�c)���B���h��*��J�����!\$�z�W/��Q-8���o�I�8&Z���'��s�zE�E��W.M�ё��S�\��j��������Z�E���s!����=����d���ˊ-�+�Vd��4���E�D��s��҃.ch�\y�Z��mp>���RE0�����D�|�������۶]S���T�����O�l���F�%>�S��r��5g?I�b��Z�� c��7��.�Scx����k�'nm�;Z��4��r�LX2[6�:+�_��r��d�g��t#:M�Σӈ�n��i�X&�ۘ�^L��1}��@X�d��;O��ua8��P�L"�/w��j�nN��� ,
Ɇ���s}�������c'����D�q������i��p^�N����r�2���$�
��q[@3*���.,�Txhp-���O�T���`�&"��g����?��1c����ꥌ�y$�N.�n$7�%�}�^��q���( ���<;Ґ�Vݢ&���VPW�(n��@�I�0����Ҽ�n�$r���u�����0�Z������x6�8�QH'u�8Sdw/�i9�k��T8+) �W�-4"��L�#\ͺ�����po���� �D<r����*����+�+F�yoa�)7�$�(j,�yBnq�\@c�}��Ǭ�CzW���	Q���0� �׹�cN�k:}W.y'%
̀^ML@�������Xke"X����`�ҍ_U�;�Q�!j)7ҏ��ƷR���M�;M����O���]�+��UME��j? 9E3Lj®bbu�$��$tT�~����ZK�5]�\��E�@7�� 屮W��
��V��LJ�B�DFŨ�f��kB]���#�J�*�h��F�TQ��s�f���;GkШΚa�I�cbp�\��8��S��:䲸�?������J]���e�$)���KK�<�à�����0O�
����5U�u-��y�Ȥ��x��C��h�N��j��q �1,�R,,JP	>��Э��
oJ���!nL�dbQ���̿$�,�e'�\Ay(�]���y�{>[@��n�d�e��y��C8���� �H:V;��eWqՊz�	���R�p'p�Mw%%L�F%�#)V�W"iqm�HP+�qKFҞg%�]XW�?�<S���BN��VX�t���_)opu5�3��Z_I�ќ[�w��:�r�OM۽�[��NzO3+�<�z2��9��">��{x͵���/��M�<��]�:g��ȗ;	�8�����s�wnkou���� ���*;��.���J���Dy�#s������j�H*��,��	��(	��2�VnOw ��}>bZ���>���wn�񵰁�(�8�OZ��D����1H���7s�4x�d#��k�����13���-��S�T�7GFC��
m�ţ��t$eo/��<�U;%��k������酵�'m�&���5�kR;Ky��`�ۚ"i�=:>+9 -!��
/����}�W?�s&��`P��x�H	���w[<*Oږ�Q���M5"o��S��^���0L�j��Ϫ4KW����X��!p��j&�X-���HSz,m���u�l����vpT�K�p�]eE�H��׀����ФS���M�\�{�k�gs��RNp��r]�*�Ξ�s�j� �x�����,lx����N�ly��~�^O�F���'������.BQsj��+��G��!��m��ԍ�#��c�� �E�����Y��/.���j��;�˕��W\��*���F��u�y>����=�0��^�{߾���0azX>��^s�6�1�l�P��w��*�e����D��|rd��t�T�9&L[�5���We�'�eف���P���6��'Rwl�#��w(i$��#@���ݛ_��_Աx�F k��"9�V���;�{Wv�������Mu����|�U�k=,'e��(C~�&�3�X
��)K�8��� x�A�qI�C��.��O{u���W�5m�����f���h��3R\v76�8[�ƍ��@k�}���ɒ�O�X��a������|�A04Ψ�{��O�'+aH�� O�ʤ����a�K�6H�o�	�=@�����L$o�gjt�4iR��S8\�2A�1c72�Z8��Q۾rô���2�w���!�r��r�i�\Fkѕ	��9���y�!b�;r�J�_(�����/ji���".ڌc�:R?��9�cώ��n���=x��������2D���%��_A�5`���R���,b�fck%�{�;�͡S�k!E�Mn�q�.�lʋ\
�f� <)�,T=�}���D���^q&j��3ɘhI���u����}��J�2��fr��?���	mF��h��#�%Z��ޛ蝼�Hm�)���޼�M��wJJ����X��jJ`�CT��_� �M��v�疿���#.�4�ЬX����ʮ�:^��r3��U�o�����\�$��5�&���4�LO�ſ�s۱�ۭ�%��EI�+�q��L=��Ж�x������{
,\Iz��f|����D�7޴okt��[q(�+wAB������[�2�F�V��fґ�w^m�?tκ��n<LT�X#�x���5$��i�����v}��4wgT":{��~�5���8��� e��c�Z4�#��i=zw3L��y.�L�wwU������%"k�e�߂`�ñ?�h�'n�P��y�;B%$�F�V��R���O�1���%�Xz��n�Sx���l�siokb��7~n�*��(*Hb:
Kd^�<q�ՙ���ϭ�3��g{b��G�εD쎻$�)D����NS:���2�jo���[��N���H����S��ogL倖N�J�Q�~�B�ǖN@dl�p�§|�S,x��cw��El:#�ߋ�=�vV�9�Pyz��<�G!Z�o�:)[��YBs{µ��F+���_D�~��=^~<��yt�w^�r�����$~VEy�kx��L��J�5��}5�{.b�])d�ω�"j)^�L�{��nF��yU���(�:ׅ�YKXמ�d�6�t��;x��?{�Y�5�6��o?W<Y��Z�!���� ��Y�B�Q�-O�p��~��u�~1�I�hz����}A�CL�AӢ10^Q<8�>��+�ZS)�N߫��X��﵌��3�����̃��<�Ń����ݖ(����{�?�,`����'>���	XQ⍀��d��a�A�E>�\Mz&�z>���{M�g/�!�W��\\�=���Pz�/��M1�W�8� ���)��d��I��bfROr�ф�91t����a�H��77�2�u'3~7CvV�z9}�mk�@�!�s���#����4��s^;d9l/l�nL�Fa���:pZ�+��,_d�N8�Q�y�z�i9�1�l�D�Db��㐽�(@�4̔����x��L>.�v|&´S����z��¡^�,C�=V���@�`��.�����la$Ȃio�%@�|$���9�.9��X��E	ݢ
/�_R��1E�Ӊ�t�?��9�D�'�R�6�F��TBrU|�s�-I��+�s������G׹�@J�zh�8D'뮇����A������i'��oAD�T��Z���w��Y	����!��w��3���=����74�V�#�ƪF�>�iI�1?0v�p/�&,�e���\�
�sc2�Jͨ�2.�P�K�&Z� !]����Y��;�39��x�l��Y�f-�AlYf(l&��M��Y�E�^�����@,/Q�3�O~y�푷$��I/�9�
�kOCN��j�ݣ��u��cN���I6�l�����M?�WJ�&ȵ�#Y�f�V�?ը�����۸�z�v)yJ�u���	��jS�1@Y�����������`0��[��Y�����<�������"�&8�[�F��w��ή�KUh>��B�m-z�t����@��S�}�M:]���%5!k35t�|����=HO�%S�:W{>T�M��������s�Ιl(3������ b9;В��ߪp*�M%U|W$oW�Y��y�����c\`�r:���9�0�~b��c�1F(������q�i�M��� P_l�v!:��=�r�>ڿ����o#2��U�v?�]�rַ��.��� i&������!L:�
���Pk�P���/*#4x}���C4�z^�A�VCS�M(c�gupM4&�t�$sbd��Gm~�sw�����/n�-s�=�F�������X�
S �VE�����lp+P���M��Zml� I����Z��8/��
J��Bх>�sd� |?����o=R�o7�0L©����=���B�r��]�$d&���ܐqUm�LĤc4>�o�OK�X?z�L����h��Ga���#�&��;TG˼4;E�S\k_�jO�f ��|ѾJ����f�T�1�̷9�i*�p	5Z%���i��
+Ь��+:�7����/��D4I�[���S����Q���ZcGY�愍C.Q*Y���V����;T'���c[�"&�e��9>Z���I��8ԘQ(�뗃�6��0�-
pJ�D�S�xw�JK� ����9R���jf�ax� /��bS��������O����k_����'c}N�G(<�^�nT�~�9f�S;���t��3�P�>���g�+o��y@��%�;�@��I�r���o�����X�!�bK����\���1c-Osq��$u�H�G���)ꭨ'���^��&�:7�og��*u�2�Q�*Q���g>����fY,��1h�Ys�<E�N�Q��L�e��ֈG�f��p�j��}Q?Bc,]�T�$=�Jm�9���.=�������*s�O��T�ܸZ��eHu�˜��B���u�_w4t[r{��G�%��P�O����_4q��u�{ҳFe�<�b�Ӛ��\vHV&n�)����$�plw� �Do�n�x��1�t�(n��)=)��bc�+�D;�)���ل�F�HѭZoU�o�$�u:F9%0BF�ZY<�ƞ̬�����.���a��ۀǞw���a�T���}eQ0�J�C!|H���K�S�]�D��C�#�ۍw���ڄ�iTL�?Cy���/��v9H� zz�\��1ѩ�$�dƘȠ�O�g���%%��++��t]r�p�����D�Ǖ,�R�{B�g!�ǘ&N%N�O#��{��g�N(K�� ܨ<Y�e��p���RY_�-�p���@���V�{UO�p��ou.� :O��N�e����H8!��g��A���z���h��ģ��2�x�U� �6�/�é�D��\'}�r�=�v����
a+�F�?���)Ᶎ��p�9�<����em���0l7��H/Z�D��V
ق���L��뛼��{|�P���~��;���g�f��&e#sD�o�1�PKYMa�f-�y]�Wk+d8+N���6ԘKt����YƜ�
��:�auzH�
��XTdf��:�.��C݇,��^Qr�33�Y`��}1�ߵ�֤a"��H?��;R"������5��ѕVF�T�ǫ	���c4�Yp�8��R��u���Z�ѐ�a:�B$A�.��5��	��]���sד^}�N�/��5/Q��Yzl ǩ�;�[i$��3|*��Ě�А�;Ѥ��гU�.�е}�����r���W��;�=�v冩�ݹ�;�}��6��?�T ����8�7�$���Q�9:�/��!y�XCVq�ËghѢޢ��Ӧ܅�Cۉ�#�A/ t(���FSu��(*���Se8����w�kb�� ѷ����ͮ��_�Y% �i��iW
\f�/3|-��D_�"g��z2�1�_t�+#�څ>��;���TR�����o��1�.�

p�ú,+W6=��!ݬz��*E`{`'�!p�󽰧>���U�Ft%�J"�.j;̭չX&�bZ�kg�_�WB��٩��WQ��!
�������ذr�یR��zY�,�Un���1�Z4t���P'�
-|/�"�"�x�����G�a9.s8�z�zڲ���"���R�^U£��ε�"���$yux�6~@�|<ۿ�X����Nw�l!�!�'�T��-D��b�"$kb(-ވ�,�t�V>~16��V�������A��(��	/��l�'E�E�Z�1���d˗(�̖nw�KJ,�lke`2<��a�6�'3�s��l�z�>����Τ%�Լ��wzL��У���+qW�ڲ'�}
8�D^u��DuP��=v̖9�����ȶ�z��� �Ժ=���w�\[5�ϗ"�i,�&��bm�8^����[�@KB����͋/9;ԥ�6g��yi�vG�M8}O>�\��ᦩ�S���W���g��,c ��ƿ#�Hse����9��H�KlF�sm�促.qYVQ�Dio�'� ��71�^�e��gD��N�>T��g�z���ǜ� �*4�<�Ѿ���Q�U�a(���tԧ@����C�|�&���kڙ9�� ϕr���q^ך@q��3�L���_�DD�-jn?�W��E�]T0j�Q�?,�uv�
}N�es�:��EBw ��7�T���'W��+}�ў�ihy)uї��h��>�p��Ek��U��M)x􏰯�%�C#HA~eG�1����G�`;~�c�kU�
�W�%���D�g��4Q�V������c��� ��GZC�&~O��MX���Q+��D��U� ����E�d�C�@���
��-�+� �Q�����I����x5��/sD8����7�?�l�K��� �y��:��lҹZ#��Bo���y������GQ��l������?������*�"E���-��n�J6�F������r,{�t��e���k�
��yl,�h�:?���!�p��8"�)�6R�v�!o�Z��p�[?��ot���D�yo�?���Vs����-`Yl!B���4���3�0躔�p�� �b���b�R��U@x@<�	ㅌ��/���(*��9�6a:��Y�է���V\3R0��)�&��L�}No�������	���j��U�1�r�Ù��H/���G����s�¢z�!��8>dn�|�����0c�+�w��2���u�����]WO�,tW���,�VY/˕�����/�?к�^�/������3@�x�Cw��m�?CT9�H�p4�]ݳ��k5�ѭ^|)� ��~r��x��y��9�M�����_Y,y���G<塽0w� ����۠�![3ϼ�C۰uB��#������<���e'��e4j�u.O��m���H_��߱�2y��f�z��y$~}0��%�]$ڱ��B��uB	���])��O�ω�؆@c��z��i��κ� D�.���)�7�K���p���Tzu��V�94�X�����>4xK�b�[fи�eٚ�iI���(\�EpRСnB%W� �ʾ,Q2�k��+�b1�:�
�lژ;�t&���!Po�,����:��{L�?��T��.���?��!�}Йz=��+;�'�1r$�t�E�'Ou�gL(���8�7�s���}�q<�l�����k���+��t
��{����_��O@�s|�c���m�Y��n����������� ��ZK<�`s�yq
K}1������&j�\v���A�f�������'y:�����(ͤ\uq��o���R�z=&7'+�ʒ�%Й��we
t��#��:��z=�ܪ��lD�x}��Y`s=h��g�j�f�)����-�J��Y�v&"X	{l� �T_��@��쟍�޶��D��� �I4�"!+�Nq�-ة�
��}��3u]m��2�>�w�+�l''�lL!����;�CEЦ�3Lj�9�)���"A�6� $4z�1X\����Z��<�4�{M�ZGH�DL� �X]�}��%��U�yfP��M_{'ބ����a��|9&c�iİz�������+`)����1�+X�
�=�m��Ԝ,�>���G-7d}h�;���$z6��J�z,��5��i����U�\��3o1u	榠�"b���t��/�J�'��\�������"ʋ�j��PLHp�D\�VL���ghQ��Y�l�������`��ZѤc��&@�/h`��G:y�ʷ'q��J�S�:�������Qu~�3�l�q�ݢQJ�C�emkĸ���������w`k��3�Y�$l4�;%�󧞓,.��;�����4El�tzWY�T�v���G�6P�W���F����]٭���T2�Za�� f�py�i놊� �0�\;vb^�	66�{��}LE)��dҩQ�YRXb�
�SZ��n(���8o#3O�Dn��I0^���_�t4Ӟ�����AaR�6y`���!G�#Bv���!i�jSY���S�"A������4���p���*�)�4�)�[w!1��z��:;����P۳ �%Ya�����M��y۰��i�c��#v�GE�$�h�D`ѓ0j����A�횺�>5���*"�� wD	���M�Qw/^�y���[ =n���l��N&����aߟf��o�L�����@��|:������Q%�+�@��T��A���y�˝�n'�`����6��L[�O�z �{}_�*Oh�қ��Oc/ȥ x��1d�#kyc�#?њ�8h�U|�.r]�ݞT�[M՘�b� <>�i�6$�~���s�3��<}��R� ��{�(��-�Ǭ|�+=�_11M	h�Q���������f�!g9&��Y����2[P��Q�yG+,$e@�A��Gi@��_w���#g5 ��l℣�q�ADx�e���4�ˀ�i�N���ǚ(,�Q���v�Ew��@ ���hY�9�R���!����=r�m)�5���t�����t'=��ʰ�Z+�iN��&����ǅ�	�=d��ic��+pw@�iܧ��dmі���%���W7s H<�Λs�Af8@�$|/��I%�t�p�p�߇�y�q�H3mPJ�Rn�x!e%�Z<�6��r�H�/���(<Y�,�R�����	���<g�ZQ(|��]��!�x���ueԗ�ƃ�-ᕖ�4�>}�eg���Ӌt��M�d������}M��S�7@��	[G�G �_�(T:~�;�f_��r������%OGOi����=��f�u�����uɌ~H(�;8;lB&�:Ù@H�.�dх�Z��&{1��y�"C�(��Fq��6������f9�����e�͹[��ĝ���F��!��g�C9
'4�hK�Ƚ&���*vK����x�E��7p���؃�)����Kx{HHThH.�d�&&g3�8_؁1����Y�4�FR�/���Z�r�2e�z�4se:7���Ԋ)�#:���-Ϥ�-�5o��ר��0Mq������l���~A��Z���ƼQɝd�=���=n�r�g��{�'A��];�j��7�<��LAԸ��
Qu'��	4�:��+;�	p���G�I#����lf[m`w��uS���a�+Q?�����&}�i�}�A�E���V�<B�:�)��R+�n�	]h��D�*z?����`ݾ����^]���{�zF���X��֘��X�-�F��DOC��'k0�$0�hX��r�����>}h��]�	c��%�NP�S,���%�rJ�JO��&�p�gr1"��3��d*��.�&��d�J?ОQ�b��\�����;�{g*n��i�W���<�c�Rٻ*t�CS�B���x�~��N��+c�S�b�zfS\�q8�!�i�CH���u� �u1��9�G
��RN�����&M}���޼�_��/gc�O�PV�gS�/�@�)�z�3k��%.��[*LC7�y&"!ξ�T��
�WG��7QgB�� �����dLTZ��ܑ �]�K5�2P�"��R2� ��xb��;NP'\;>���[�i:0�������X���(�y*��F6���<bS�,�C4>��Ӌ0v\�`zq�hY���.�_��:��[����:��U�c��k;�w�-��C�Mr��rts����
r���e��q�?R� U���6�����+�1Z瑂��6���kh/�ۭeH��K�'�pR,?.�I��>��Z/��Ys��(�R��XoA����\��q{O��b��	�����<�M�VGt��L>v��])}Gc��Û6?`�y�Qм��c"}c�����=�pN���E�]�;w��;�P�)%��*����ĚNt�a�W.^��Dԗ6��������Z(�r�NqX}���ܸs5��~{Y����(���y��e���,���u�62��7wz�J򘹌�5�p�4'�r�p#8Cܴĸ�����hf�c����"����v�0=��P�����ƣ㌝�Sh�7�Ɣ�N�~)ia����T�O`"$�L`�E��9��{�r|k��g�bD�/�[�~��{����3YU@�Q�/?�ᤲH�73�pj��l�r� ��EIf�p�t���'��{,L
TI򿁉\�G�#֐����)��Xy���`}a�c�;q\3$��䞃E����9;��L���aX�6�����B����Uݽ��#`(N��+u��%hm�0�3(�j'!�P28-��9<<w����n��̧�S��*ƃ$� �;Wlȋ>�鷸��έ��K��K��