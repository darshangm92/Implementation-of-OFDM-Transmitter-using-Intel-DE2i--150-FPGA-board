��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<����貖���\&�
9ڠ�D���J[�J�\bT��0�o�o�o$�t�3�A9 e��q��}�&����/	�{"'���
��C��E��;��ν6���{7��q���Q�JU�Oz���!���5���
d�@�1)l�})��X
Nz-�&�=i�R��,/l��x���*Ɯ�{�����[S���Ԟ�{S�F|��z�,B�<�~���Uߠ�V"S��eL{{?���2;��l��`�;���p����|	�����U��=��Þ�����{P&�EF��rP�l1zoˑ8>�A�����E�+f�"M{���C���2߿�ʙ(�|��r=�M�Lز�6��jo]Z9�V�WA(��������Gꉩv$�
�?�./�����X�ʭ'^�`珄�4�õ�~�%�z��)R�C����\�W�͚B�>���!zі.��Αe=L���2�1����� ˽
��J��"�.��)�&w���+�3�K����vG��H��7v(����_L��f3T����4-֪^�S�b}���/8#`��b�m��䝑��Tu[V�vs�o�]E��
�,�Y����a 6E�U=s5�!�S^u&�ϡ��� � ���%�$��pΣM� k?�-�Ge�����M5a�u�2��}���yٗQ�mR��,�r3�l�!�+>彞��3>E��6��RN����ݦ=j�N��y-;�!����)��T��q�E�Ale���&�HY��Q��T{���i�dL���p���W����2��!���o~72��B`̲���ԇ�ll%��EԗC�X���Q*E�HC���S16�&������\9P�*���"��hZB����#?a��U�O�>qw'���.:6���Xy���7Z�-Y,:�A�I���r��J�aF�?g]Y �kQ����v���g��&�Pt�3���-��M�4P:~���VG��%��G�Q���zՀ�VaB��o�%�w�qÌcݱh������>�!K�
�#�5\R�2��Rf1=a�\BF����Xn�m{�G��E �It�&2s-�O�	����N]z'��J����0_���h5�Y�7�?��cS>��>s�ݷ�;&��vD�h<[\ӟ��Z?�y"{P��`���S�eA�%�j��_Vbٹ)��K�wRɛ�����sb��L��r��YB�L\�AR�����H�����}�qNƦ��Ͷ�P
|dϺ�&c��y�3v�3�F���Q�}�zI��!���4ʥ&��Ɛ/���v�^��k�G�������7�k^��s���
�!�{�-cr��*P���i�B綅�+�B�.�����$y���F�ʹYA�?�F��D�Y"��fc=}�<l�HL�?����@T��,���x��$�y3.��;[n��lc�=������Y*О`�o��s%�K+orP)f�������Ri�!�X�!B�V�h�#�������9�2�?��8^T��p��� ��hxk�����K���T���pS��fє�~��G���"��d��y����Y�Hs�^V�c�4�Js�j��L@��f�9cރ5U��
�ʵ�Eze�r�n��u���O���qV�kk��ϑ@�<�yb^F;��Hsi���Q��������kM��[��m1��B�-u�zi��dg��}������(����G�ߠ C�*M��l��:b�����N��C,�����O�ݶ���WJ
���d�]�y�t?!�Cc�7���P:��\�ll�H��T�l����´R����г��~���VO�N)KL�{�vLn M�/�X�lG���E�T���L%tt�̭���]�|.!I�/.�sF9����u��Ե��kq��^ąe�7�2�;�c��D�U*�%[,�z��ПN�8�x���Rt�}���r��f�E }3�P��=Xv��C�e��๳Ou��	N�^�!�rA�Б枅.SAV�����p:"2�jj�jl�^�^���p^��>�Xg�(]>ᯃ���&�c�Jl��.?!w�e�\i��QC�Ɛ>٠i��
Z���`�+|~�,W�f2�^�X!t�uг�s�¸�c�=}�#��}Z��xSB��D}=�ܶ�ɀ;�o�r�A��	
��|u��m'���u�`b^�Qq 9�����ו������ץ��sC����^��X�Qm���c�&3j�.Mߚ��T�Kf1Qō]�J�#zG�w٤S�t���dq�J/:D�9��VQiSjKX��{����U���9	���V�:g��cxj74q�f�?��*�}�������5/�+�r�t�pU��v����O���
�-���*��� qG���1(�Nٖ�t��2����B��T����7k5тo���=������)b�B�L�v��zS�{mx3��^����͋��7��|~�Gb��¶W��)��jq`�(v	�d]6�=[���u�D!d��o�?�l�d�6v�^�Y4��[�49LD���D_ ���H�b)xv�n��%[��?�`#ҝ:���ˣ�����I���z���)���M�6�.C{
C���޸1�t�>vs{/�NZ�p����D<�������2�Z/f���,�}��7S�=�+��@l��Lԃ����PM3�u՞0<+�Lqܕ���-�h��.!�p�
ӭ���g�݀���N�]���y�r�|k�x�|�5������r�Ƴ�ÆYp��3���o+������8�:˚
��]z�����v����+7�`r�}&�>�"��r��O/[�~%�9*��YP����H�������uՑ��3l8� D�tS����h���t?����x%!��X5�f��L�����Y�AIh��Mü;��G��Æ��V�%�V�1*��gL@9��u1:��=�%e`Z���]Pj�5�9������~y�
�uP������u���
�U}�I���zbK�������?�¿�[�p���W��-_Yd�
	����
��m�����>@x�5�T8�����$-�����l�n�u��8�I��)l��KvD�����zL���gr�-Sj��m�51Ql����ux�����E��>���B���������ب7��hvmz���;?�0�$ͽ�/���Q&�����t\��㖨�l��n�KV�p\֋Zo��.ļ���K���t�mD�q(���V7ʽ#���h���k�HM!d�l�4���L4��9�w�I�yE�uv��]��g>K?��z��R��x�3�P&`�:�'��$�$2���Dx��'돥�^8�ğ��~�^��C���>��Q|����:
,����$E��^ҳ�;f����_�s�"�r��(�Y���>~
#���P�9݋��ED�j�@�ȫn1ƕ`7�c�>�ǎ9 VG2�1���YG��A��M�&<�^:�>���otPj�$f�}HdJޮћ'��s�+�h" S�0�Nv���ί6�F������z�k��������s�,�(�m/�𦉨\�a&*	��&P-��j͏3.�%S{�Hj�G��>��v҅����0��~[�%�C�L���Ƅ5Xv�7�9P[��^��\i�������7�M4v��1&G��$I^79�cB�#A�J��U��g��-�?E
�a����z�W�e��8��|�o~_XR����$A�"�*���O�Eru��������Tg�9(�(G���|�N1� /_�V}d���;��	�Dq�x��C��������$��0l'��QGJ��ԫ7&�d����K�\J �{`5�˨9b'7���H�����/!��*b�t��b��*���峙����Ο���R���Ab`�t�i4���>�Z^I�R�v�4D�26k�5���J��ݑYO)�-|�#g�a�^���^�w�d����$de�[/=ũ뗡��J���8��	фw濍�_�xC�z��D�N֛i!'���o�6KNQ�ֶ���5OsiB��\3�ӳ�,mw�~~��y�E*�,��|슶���
$V����,��Hh���Z���X��'PM��"Ԛ#�A�(}��+�ޅ��Pt� 3J�	��i|�NN� h\|�B(���K�:���)��Dy;�rgH��f^
hT󁷍��7;�mv"a��E�τ1wu��w'B",2�Cl�k�t;�m��z�=�'�<:J<�� �j�G�h��U� �g��C��P��ȵ�����{��ӥ���F�&��h�p: ׇ�l��v�Y�j�3'��N��F�T�#�y�K��ń����<2���B҉� v�Pr�+?B�('@OQ��HZ��Ώ���"q}�]L��=�e��(��(#�uvG��ˑ*���~$������ޢ��*l�g�%�tc���,)&�?9ẩ���D=c�����*�jp���l%4����8�Ѣ]��U��j���[�=���4����z�8D��wPO�%9m@�Q�-�<�4E��L�ވB�!����ט���>�� �tqƩDN[�$5f\\�uZhtZ��ƴlV�kjЁZ������"�S"R��K�Ҿdb����]�ϕ0&Wyy�YA�R2|A(�ݰ7��F�n�1����?��=����<l�� �V�h.�C�p�[���R�w���B[�U滄z���.������(Nh���)�!�z���c{P���� �Dg}4���\��;���.C���(k�o��
�X���~(���L:���ɽ�$q��������o\��"`�\���=@+�OqZ�3�a
E�`1`~���#�w�6]X)�v�e
���|�<������#+ �E���,`���k?Kܘ�:�ś+$��Xp��8�����h�U�ۺ6@�T%���p�54�o�R��+x�G'�mv�wI�M�:1�.��`ԮJ�}N)�&0�J\�ݻw��,��R�}ܳ�k�BJ�"཭�t���Oi�O���V����a����L	�@�����lW�(�81�<$�f��tF���K ��x>V�@��O#mIM��[bU��5�~PGobIz��~����._��S��Ԯ�$M�_�{#O�i�ȸ��FD�q�b2����d2�cP����n&$�2����cQ��q�q�����OzN���V����9rĸ�ܜ �h�����e�����������ƭQ��J�K�G^)q�+�g^������\����O 8���_(�9F)@���K�J�q�e���H��gu�C�`i�g��5[yza/�8C33uO��kB5CJHB�&7�MU^��~_5N��p�RB��QA	�+�weL�4�_Bm!<Nx�õ��6k��і�D)jf'?�
�:axH����M�}�[��"yK��hwt������{�v|0���o��5��}�oi�(QF�S�U��]c�����\���is��k~�EO���xi3� �O9��w�:���G'�Cb��r���6}�,��(U�1���c���z���J '�@��ޭ��������VU	��D����)io������"C���bۅEB�Y�r��Y��H`}Ão��r�[�
k2P���sd[ƮC��ѳqD�k$y�����}l�Q�q����k���E�1>��M���A�]^Ȳ��)�$m)�r�O��� ��`����$���<l�������ԉ� u)FQ�?��.g��M0��Od��0�8��!�򽎝�m|�8�N��b���u�C3����c4�R�HK|���2W$S�8�衭֣�%��8i^9:�����=�؋�-n�=B��R�6����]�.S����F�<�1�/���}	).��s����c���;0�ߎ�B�r���*�.�~B�^������<�b�e�m�'[��HC䐳���$��υhr�On�Y
�O	�f&yv<b�}�<t��弿y�}/���~��=#;3�����0H4�׸9���d.8�'dtȖ����:qG�:-A�irD2�����2��he�e�YY3;���N�����s����@��dÜ�� �n�����P5�w��)��n�n�F��7{��E}Az�=�
Q�I�Ӷuj5ˏZ�f��pВ��C��鋧eb.u��VjH7��
�k�Vi����B#�>/>�3��=8���q�w��&0R9D,���fÚ$ޡ��n�� >�<,)���l�ջ�I^�����h@G��R�F�RLU8�0���i\�b��ɊI��LG)�v�,��e��wb����ڷ�%Y5 ���z�k��?L-��p�t7>j���׿H�LC�'$yг/�m�_��pq�ʟ�0�u~UŵGd\�S��9ؒ_��M�4l��+�5�C�R�LDz��+B!(VvN|�8-�5�'i]c��qw�����&k`{:X;9Y�0fZ�W�(�9e�����!Vj���F'P31�*c�^s�PX����9�74<��;�|�^8��5���xWQ)�ˣ��ޛ���-��a�����1�Ն^8��W�{'ۢ��w�?Έc[7��V��&M<�����ɇ�8���׈F@t����Ê�+"��/�U"�a�b��F�__�j�s{�d�-3ѿ��JC�w�aO4y7�ߞ�K��k,��`��L��Oh}��@��U�!�8��ǍB9X~���=-��K��>	ꎑ�uYwC'3�G���G�A�֛���uK���_�g�J2^f����kW1֑~N����I�����?R��<"��Jg�Ր6G�s�ӈo�D�1�OQ�Rn�9yS	������