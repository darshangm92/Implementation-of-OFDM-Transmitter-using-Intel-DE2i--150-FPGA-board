��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����G��՛��A����_���E��{�o�j�-�wmy�#fnqąMu�=J�(��]�
h�٤����[��wHOWeG�# ��'Y��l�ݱ_@1 N迱L<���I� �9�F3�6'kn��[��cv`�Ǐ�՝kb�v��T��mE��oTr��3a9��p�	��.�� 1���s�.�4�ra��������K�1���ݎUʐ����v���-�W@��S�'��t7��W��j?Ц��5���@��������T���goL/�`2��-�������ގc}�39��-9K���b��7�r�^1(N�o{�!0��Z��-�/�)�;���e���"��P�+r �(����s%|ǚ��
^!l��$���P�1�V4���p�$Lz�@�"o���.T[V:��W�(�q�f!�/�Β���JNTF�I�����^n��LH���QE��7d5��<߂�0,^P��K�(a2 �R���Ay�RI`�Qԙ�n�Oz�C�r�����8�Z296��k| ���1.[���$���x@w�2��ELL��7,i{��&�W�sG��gzE~K��i�B����Z�N���yf�Uo�*�V\m��)�b7�	q)��m.Hm��{ʈi�O�͇4&*�)d�6����Q�cT�J-�uW�Q-��+����B�9��K��m�c���1����'��������g�{���>n�.`Hnn��D���Ր�mK�a�*��:�l����'R���)�sf���آs�V	J��,WE�M���Բl�h?ŒZ��d�/���oW�xC;��H֐��"��J�W��0��@m��q.��<����[�i��5�{nrYl��hKpǚ��L�<�Y��W�;e>��4�m�ĤV�,L��o�A���x\��d���h�8�Z�V��@.l�A������I����C��`$Q,~	����| l��BĜh�h��[��y�e�)���t���E���k�4�6 ",%�~��9���8�y��"oO�����d��6:D�L�[h�U�Z��{'��r�,]��I�? и)���ԃ�	�p����?��1v`�z�u �2���	�#���O�G�:�1�r6(�8H��9Tou�LV�A�ϳ��,�����+�5�/h������~�wd���Y��1�(�_R�y"���s6�VN���+#h�H����II�Ȇ�������2��i@���Ӡ���J��Q�Ě�丼U9A��B{( ���ecS�L;�mΩJ���w��F�yv�	^kO�#@����6�(�fjѤ7)�.�	�2��B`'��/-v���������?8�\���֖ŤvA�:t�X��2�.i�����; 4]Q*����|C��m��I>�7XVI�"�����\z�q^&�{�K��G��J5��*-p��W�@W���NПEF\o�+#!)Y��/)}�H�y����x�9�ع,�nDI=M���ڗT�,����(�u���8�z�`]-3�F�NHb}A�;oNj�!NcĮ�>c�%^d�����p�y�HyR���~N��G�,��3���1��*�9�o2�X�C>9��\S���e���-�tؽ�#|?.�v��c�H� �Aj�%�����±��#�ayj��28���+��0����pߙ:��DV�=�a�9�C�H�f�E��*��9�	������S�mY2wUsBrxΡ�[�)YuSY�0�^#��7X�Th�w�7����N��4��v;�N�e�yKy?���L�ɀk��p��|p���{*���Vs'a�r�*áj��*��yp_�E�Ϩ�F(�n��m�ފ�1%�U:.Z�����X�(<a�H1���"	I��X�ng�q���a��}7��ㇹ�P��}nԝ� 3��m��\��0mH���� .+��.$�����ȍ��3*��9I%��V?�hB �ךR']���:/���=���ً'�G��s��x	48�)V�ٸĶ�Gg�	�/����I���?�;t±S�]���W�K�fm*�]���lV� ���r7��F�f��?q.��֡ &��ye5�mW�,�E�\�R��(�����%��rz�~7p��x��f��P��BƖ�G��C��b�~�M^�k �Vr����e����kj�K�@��Up*`��9��A���t��W����O����Y�9ے���:�͝�y�t�����2�v�д�!3%S1�l-J�/� �3�]Dz�d09L0��)'�Io�p߾���6�@I���L͟;K�ɠ������ɦW��Y9�����=�+��||����p����QHxj�q�u�4���ȓQxcY��(�����Ȩا�}V�<d_�̋k�
�(W��=�QH�аGZW�#�-ј-<E[�J��Y�3LB"��OA��g+��'�2;J����� �L��I/�"�h��:B&]!�<hc���Y���c���25٧F��;Ud�\	��V�ѧ�ƭ@Ժ��i'�@�Ƭ��w��@�|H�W2�'��Z��l*�=�SY�_Y���Bj�j"Q]<��.1ڠv3�f_�p��ҵm���T6����°(��O 5�������U��������57��f�$�-� ds�g(��������	GN+��,0�?̈���Ps@��wP��B�EY�_)�'�������v�
P��^�ȓgk�F�f�(~;d�j�Z/+�ײp�,���I?t*`�����D"�<����iO{�bDW�4Q�q�T��SZ%��l.ϧq����$^ej�j�|��$e�ͭ(����	& k�P�������/j�D���K=�1-�A�$>Y�]��g�1Z�����<S�ȌѪPa=67\h!��`ի���ڨ ��Rd��q�)�V�yJF'{�!~E��eS%�W��Jɽ=81���
���+rS����T����r�2S��&L�Zw�~�<���Ȣ����.�ʟ?i��
���hd�>�>����\M4�_����@#���0�q�p��y�Nǅ�Z�7���� ��H��_��I�_�j`M���b��2s/�Ax�HS��g-�-��b��1�zm�����~���&��Nڽ�#=o�Ĉ h�πa��]���\�-��+;'V�qX3~���+J[Q�򑕴%�A�g�iOZ��Ԗ(%g����?�F��x�z����Xb�I�V����ڃ�xG��K�2~�!�bN�X�eb���Er�TD>��h<�k([j�0�Dey0*Ӝ��\��X����l�z6���F9�uI�	֋�捯^��s����)8hkg���&�|گ~B@)udO�>	K��w�FTdӧ��NÃ�q^�T?;��+�lH����I�fM��慄�={B�os�YG��1�,�.p�X�%)O���p�	���ӕݪ��V��J�RTvՃ��m����h&�d����� l��J�&�V����R�J�m���)��L�W�
�ǷE�sL��7���e"�(l��s��P{l�j�c�k�)#��n\���&�}9��2�8�c�3�yo�)�����x>�F��V�=��+n_I5޷�3�4��x��	�	6-�B@���5�2��� +-�Z�t�(�FT-�t��2�<�,:�#��'�@�=���8b�fR��r�J�M�o�k6��Uڝc�j-�����J�c1}�q�Oޕ�u�Z��g[6��(K�����õ��k�G����V4���'�����⽁����)a���{�����68N䬘\3�:�WQs�]/��3��>?.��a�a��?�\L��
(�P^Q8c+��`���T�����^�[�h�T��(����<����E<����S[n�gL3�-��6���䩅)�"��o�l��u��4�[W�_����Xb�rɁi�l+�Dݿ��w����{:ڙ�ʿpRUM�0����C��J�D�(�-O�3���=�O�-{���Fϭ=�wF�����n9n��Bsu�Z���:4�q�t�ڤqv�Wb�5������
([ym�F@W1"�KN�����y1T�_�Ӭ�b��ݩ]��
�p�f6��H�Ų�Q��c��1��=���
2�.H<�j��&v�a"�WBT��]Q��+IS%N���* �n�m*��l��m���o���~U�AV��˝<���-=�=O�B�}P�׋�#z�{��h 
]�RZ߳�K+э��[�c8�'�N�[�E?����B�B����{�p��������DUz�)p��A"��>�L\8��tH�:�",�4%�9�%X�)BP�=�k_}szD[�ƺJ#0q\�"Uh??%��ǃN��D^�W�/_��(,����p(J��u�'sb}yA&a���S���L6���	ٸ�2��94(v�Q�Ɓt��E����>��#b�>�%�ϴ� ��� �I�MC !&c){��,�f��Dl)|��7Zx�=-
2�F�'G�M�_E=3.�ֱ	d`"���� *�t���ї� ;}t���#���7]�?�
#|��<�x�}�(߇s�36H�8kZĵ_&��{� A&�7LI��^���hL:{��/	�ִ��/�YR�+,WlP�a�$�9���HFZ=.�&�b�U�l�&;����bYS
�G�R�M6b��<r=�I�Rpj �ngҜ�������S�A�߽��+�|ϝz�p5Ƀ	�ʷ�?m#\{��EV��5��D3 ��V ��X1q�'c�J���T���D��o��.PN�)����-�=��5���	g��n/��{��Jf���� � �u����72:�jkӬ�l�����3C`�Na��x`��d�����]՗)�8g�GbJ�޹�9K\v����S�x��#�Y�d�V�3���*�r�$b�:�o��3��V�7Զ�7�1��ȿ�c�Jp1��9o>�)����h
KV�ߏ�K���"a��X5`���T�a����h��J��;���m�·�`�8w�[�:@?Eɐ6d���������/�O9�='ܽ�+P՛�}}��L# ��m>��t��"1j��y��`]�XQ���{ZP��?�@�A��	��Zb��W��9�+w�����%��{^������愧|�M��ȕ.m�Pd�⥡�ב4-�\n���Od�r<܈���V�vluE-�/ݷ�5͞g���L�Y��s�s��n�pӄ�*s�3��/��	�0�XKY�s����6�l+���@�C����Y6��Iq嫁B(2��z�2�s9�x6�3�Lͫx�X���M�ow�� ��p��v��{�Y$�mpFl�n�nW�������ϣT$�fv3~�~D��=�Iȱ�3{j�ں�)f/s	��"[��^�����=�a#�f�5-���#�X����
p��D|�q�aK�A��|zD7���0���yd�,�4.���j������tR��Z��E�ؕ�e�u1�,�9Fs�K�s��Z&��M�ϩ�a�r5&��Y�s"� ���)k����ƌ�J2Pi)���O�kZ�+Z��Qؾ���u���<����@�p �q	V�j���(�i���ӫQ�=���qCRJ�ՠ��q>� f#���f��Uj������J�)���lvt��?�^��]3��)?�����&m���F�99xZ���@�ﻵ��۠�U����a���)����A �>lׅ�|:&6��Dt&�飲7ܒt
��?bj����
�{�s���|��Ó�"#�&N��8>�7E�3���?.���-�4hN���@K�y^�}�:s��4_9��:(�,��d1o���yj��o�+���J�,�S�<����!��u`�j�U�x�~��e2�I���$?�k �0��!����u��*�"d�<pw'%��A�U�ř�+= HJ!�W�n�J5�g�
.��I0�b�ԁKBH3I-�]}�Ւ��+�IT�ߑ j�]C[֔r�d�$'o���# Mg��I^��?��6k�����<|���8p�ަ�8�d�T� A�?'����a�lm�s7_��x��T_0{��܃�GQvիrn(��50|cf��=�(��#7�\�0�<*�8�����
��9�LJj���p$�������qB�q323 b�Nt����D7�0�iu���􀟲չ�"y
,�Id�&М���"O{�����2��'�pT�R���W�����A����� ��`&����'�ה�>y�U��`�мı	���@��� {c4�����;�X�M�U.V�n鲞,�u$�2gW���Dy���odK�����~FY����'��h8�r0��R�)ͩ���C�r~av;v����"x��$7�mU�����e )�ߕ
Z<��k3�y|�w�C��N\,ua0�p�I��Pfk�p/P���˸lU^υۆu���������1�~w�r����h`e�[.�.A�jU���ǎ��U��@�M�o�8����O3��Yz�؅�Eh�h ͚�Y�&��S��3j�RL�fXOZ�`�/�5�dn&1*�wS�sU�Ǚ���w_ ~�$�����b��<�ș������؂��R`�J�aĽ�η����Qs�����]��$�(��1����:6Z��b	�)���l�}?17{2Zڰ���/q|��� �2�s�!�ě��٩�C�@��W~`�/1怞�F}_�rvsԪ���*eH���2D�V�H����&hb�F����ػ~���F�x\�oly��F��ʘ�ėy*�p���5�'O���q�+���ӓ�=\xX�����FO"��Rn�-(�K!2GS�RX��*�"o�r0�4aT�	�+�P��db��$yAj�;h"���b�#��#�/bt����V޴�g��n�d�`�1���J��,�k����'�7��ϗ���lT�y?��XC�zU'�#�nV�Ó�X���1�b����������,���� x���z�2r�����_L�Iݗ҂.
��H��E�v0�]���ai�C�Ϥ�Q϶f�]��ma	�[#��\&1-�v�*6�sǒ�5'D>X�.�)7�U���d�mw
������������S/�Ng�^��r욢�1
j�#����$�ʪ��U\q�����Lωc�!�u*IN�|/B�,�X���{��x�w��� {@��]�^%����$���9��y{��+u�
ՁՄX���=S�F^[����$���b`���?���@�>HP�,��Nk���;y	8�n�v�4Gb	ΈyuS
"2��qP�C�E������`b6��p��0�c ���R����� �N�Ρ��#H�;�F����nB_b^s�Q	,eE�`H��x��M��<���b�q��|����B߲�x�k�9��&�.�TD�y�i��at����C�,���aZo�Z%N��>ȣ����f�Q��;o��朔mO�����7 ��E�w��J�d��T�;�o&[E�6å��:=�Y�l�UE�� I�
�O�08�R
L!!�W��;�*�4���~�L�g屢�:Σ`�̒���'��4a��h��p-��C�M-Ag���4S����_������[�V4&���'OT�"��=�ޚ�e\���[	K���I��?��D�(�r��٪~	P��ot7g��H�̟n/�+���U	���.���c�kh�����p�1Gi��0�\�z��\��m��©�����y�Y+"Nı�._�{��M>�FPIP�e k�;���U6ĕ�(��wx)a�B��"���jٝ�i�ʯa�f}��y�^�ފW!�K���2��$��_]��ޖ(^q+����W����oH޲�tv�Tp���Ao�_�)�%���;4N���?���\GSd�S���y>Qv��o�}}#݇n�����;�E�H�`�h�K}��(Ne�Z.�ī.�`
h�;�t���C<��#ی��#��Q�6(�b<�G���Iٮ�.�����/ke-j�r\z������L�QFyN�k�2W�T��Sh�	ñ�܅�q��*�6�����82Fa�S^��TG|��C��?|_�)�8璵��F�ߌO��ߙ�0�h]��I8.'�C�ᖄ�'����o�D"j�T>̪Qt��ie��v���	�vy��~[n-�ö�E��5�%�%���F�i�g�!)]�`G؋0a�]�v�	Է�5�W)�����	g�)��cN�I�`ź�K�ɓ�*t1�ّt�0���aZuMh�]���m �3)BkՑ��.J�߲�M>m7o����3��wp�VR.���t�;�`J������vwdhG	��7q<fh��_�\g\�p;ys1{�V��ϷT�>Ք��É�Q,�t<��� E�����	ۤ�Oyk<,<I��c0�y�'篧�ļ˨,��H� w�,����4��+��@�d�[t�U� X�[ �`�}M�I�Gn�4��w~LTql��z�޽�ġ�ϒ�u�K����C�c�͡��Do���g��f��t>:B�'��q\StP�Z�4O۱N6�ޞ��|�O:��hƀ�����1(� �����D��<C����g[9D�ḫ/ �Aڕ�iH��i��:���M���O����~�Zޕ�ɭ(/�m��AJ�D�u�Um�+��.��3���|���|?�l����!�q/%+(1B�S�?��=�8�4h�~�,)\\I�3X�y;��R�!\���m�L&�33�%/���T�J#oFS�e�Vy�r=�e� 6���eDG��c4����\�|\�:ݺ��ʇ�D��o�+}�:�h�����#[��"M>A����Q��sY� D�/N�!\���O���)��[^��O�W������"�0����n�O�8�i�!'9��)7����/�]�U/������)�$��24��)�;����΍6>���6z3��E�Yi#��Θkg�k��N\yBE��� ,XG�।���hެ�$/��M��r ��-}Vy���uSt�T ���=U$����W�`l��എ��)�R���U�L�S���u�X�眬���a���6��F�`�r���e^q��{R��N��Z�0�t1C!K�SK�X�	г�]�n�����HiW��$�P膕��:���Rh��jS�<g�l*�&��̽�0kűHx��]��Ǉ���2~�]�O��`8��s���������X�s3�6�F^��0h�R���V�k<��q%���Wl����pZ�l9 j��X�	�;-r
�<����B��k�Ej���&����jgE�u���h�����߲����Vʜ�!¹vܜ����6��d��,�;���|����Fxϵ�JZ�*�����v��dG�:��1�,�3�������&HԼ�pNv�ms���>�#�Q(h�����S����_��du�uoИ&F1K�ծ!n��~������������_�����j�gd�i,�� D�"^�&-"�$m� �W��c
����OHi*v�W ���t����&#a��'����ٛb������G:�s���uBsZ�w���0싸�e����(���~E��xH:�[}4^Ο����'��_���@��x���o�1��"���l�P�^��ږx+�4��2�0�XE�Pw���<�"l���n����%�'�Z����d1�""�!��=�-9��
|���5���t�+3Ma��9�r<fzJ�t ]�]�_��yW� +_?h����X�?����*K:������9%%�Ș�mJ�����{��z�vX������h˩F5(�~ZM�r��b��P �w�nhSzq�M2d�O-H�bS�������
��xʒ�)儰���8�IG�m��J���;�)�̰��P��n�2��!�}5k�*�ʼ�b"��*�XlMKE�?I[�}ną��_FG<���K�_�_�)�#�zP"����$�~� �T�n��B>��|lm�00�]�v���8obo�$��mE,)��"֌����2W� <�0X�X��u��{��0QS���K��m� @��9#"'���u����2Pt��d�w+�8���1� ��e�OA#�!!��Qn���2� ��\�����*�|O1�jN��;J�Tl�Mm���G �מ��A�L&-��_$��q�Y�	��c���#0��տ�ܞϥX/�5��>��=��T���!Т������@���&���m��x���;x��<3:��nI�uge8܅Ï�#�~���D���Ց����l|�2}��%.����.�:\���S�i�{D�O}�v,�~>�r@������tUYn��S�KCL�s,���;��:V���J!�}yF��S�A�۷�0��6�:����foaE��Jrz�`杚<�D�o̹R�g��[����
�q�:�����V�:��lre;�0V�S��o�+Ajv�U��D'PJC�V`�D*'X�eez�a|�3��#� �QiO�,���9R�jHa�qk]�on	�M�У^�e��V��q������'�.���ۘ��]��,��%o!_4�Ķ|�XYVʷ���"�}�S�S����ٹ�5��	6YwH�ؒ`��O�I���G[��P�k���G�8��i[F|�U#���@������n��ġ\{����8��5��~�Ν�$	C���XۅRO}�wa�� �������ix�Y�6*�3��.1���|�G�Yܙ��bs�Lk�3Gg@�
KG���VM�>�&�O�$���D���CZ�.xQ�tX5܉<:k�W�i���t�j�����Z���̗n(���I��}j�?���L�����;��7������Z�׳�f=�`ZFv���q�#�ޗ�y>E.�����Y��d�`�*�&��~�,*�-�v��a%����,�J��!�
�iI�Ǭ%p���F�aUT;��6T}�	��H��]�ݏ��\���״<ϒ)�	�S����I����s�/n���ud��Ǚ��-ʠ��>y��(q�WSL��=*%'��mu�Q�k�0CVVe��B�ʯ=���v�-��8���%%^=t����uW�����M�aa�f�@�����;CN�S+����T�K$�H�d�7	�')"X̗R���E-�֝�*��m�W�A�%K�6瞟�����Ԣ� ˩�܋ՐE7qߨ��zF
����w&���5�]ȏg
f_Rj���!|�\�ZL����,}r�#s��P�~�B��<BA��K�v�����h���*�.�aH7�	��ܿ�1 ���Ύ���~~X;�ީ��?0�1�J�~��thKu5��2�gS[f�+~$��Z:Q���~L���OwY/�k2�xC�M�����*`0#�n��2b#�Q���	����~�����P{��� ׿��h8�v�.Ts�g�uHU%��m �qm7�����A:�4�H��X?���Wiu.��P��$��ɽɺZ�R��gPU͞�lPVK�s��a��y����$�4��@ ���n��/"pF"e��k��m��S�Z��:��4�jr�R�5�ţ�d�(nAB^y� �
���,�ëٷ�:+�K���[:<P��F(�#�ş�s1)lL��pkDH�=&���H�x����;�QߘxĶ;c���t˼����~}�[wN3����[��=.Z������4����'�����[�7�P�+������w�Z��V�6��{!�Od݈���zB�41�d�8�u��J�K̛�췃��B0��>����%
q�bt�7M�o�}9�k�kpU&�G_�������Zs�轸
��T�T���T�h~�ca�aQ�۠4 b��=������J�c���y ��{�ڢ�j�Z�`$�I�-}��^S"�"Z.5�*2{���dV]	�ǝ��0$g�H����{��I��P\�a*��Z��<���j��9�C<w�L��a�a�k�A�o�Q��1Y(�����f�`y�J����}]��Q�"�}�l�<-o����	��]�w�4�w�">��L�أ	�q���hF�#ܳ<.&ݓ3�J��d���k��.�*?���8ާ�{̎"��QQ�DN�!�h�W?��\r�������X�
p��ﳠ�"j507�^�*�[C� ��'Qf��[��τ�����\=�ǉ;�΄������iǁ8QIf�VyŸߏ���)��nZa�����_���- �מ�_�R9�]v+�wa/^��t��>��q,d�K�?�F�ms߼y�`}��A�2��<h�<��?SKX�T���{�B����n�>V�1�#V�o-�ܲ(�븴`���.I�o�ƾ�4�&Mk��G�+T��h~H��;�A蒘�x��z4�('�R��`�T�)���(����<�� <�� ���]UC��y���#�[�̱���M��E7UW[��Gy}S�$�����	bX{�4 �Dd�O(l��FR$?t���|���7�M\��}�W�7+��ˮ�HV�Ptgh���<���ӑ����f�B��J���t��I.�0YDU �ԗ7Kx����-%�^rb%dw'J#����p\یM�}���+*�9{��(���g�L<`n�\�x �,������Kc�T�m���T�Kl�z[����S�C��a��N��ˢN��MpTGj[e�/�&+:�#1D��%�������b�z����nBG;�����������螄[�'J���6G��F�����)��3���ē����`���_��8�������zB}~�X��`�G�\��P������m-3�xI�G�Mx�z��c������]�ۡ��	���h�I��;��;hʕ~��(��}�vl��F{��������;����o�b�3��'=��޽�{�����tͽ���1��2J7�h� �9y_�84��acne��MCF�>�s�t�-u6�9���������p$z���M����@Fdo=+o��&{�t�NH�?��~=���\�����o_��B�|�;��E�]�\(�� ���:Bu�/6����k�[&�4� L�	{��m��7S�N����ˊ�uGb/*`�c����U�w���R��_�H~C^�@��Jۨ7.���{�l��"��>����tc�nL�
Ԡw�����k-�g��tά��bP夫��W���W����O.�[����'q CQ��n��ym���.��2P�x�.R�fg���������{��i���U�����29<����C��s�yُ���nT��'�6���O�5+��b��� {1c�(�WVx+�@BHt����}R�^oI<��񎻮H<���0����������g�u�S��'��^���G0׭F� 7i:��>��)�����>�ǑS�K�|\�2�̄#`@a��慣�� �}/�����~�+�Va+��M�}��s�+>���p�)���I�oz]�Yґ�L���B ���c�`�x����ĚBN�`�xRx�B�Y�;��)0��2��L
����c�l�$��k��T5� �3�s�of���������W@JBcL@�ǆ��g���2��y�vY�22�����Ļy��e�7oN}&b�zIH� "Vi�?%�5�n.- ��)���4X�����5�Qc��_�gdϰP��2��%������wȐ��mh����޲_rA)O6�|ny;�5��S�n�R�S�|��1k��U�R�L����&C�K�3��s{N�G��mz�e��#�N�zӾ�&��ǭ����g�%�A��г�����P����r��$�#a�Bҳ#�Tˏ�x
��U5T����˯d���.��s:���ʦ�n_� ��/cZG�z��F��)�5t�%$D�(�;#�NM��y!cD%�$KVA�@;)"�fK�A�<�<4U�.sJ�VKvҠ�0J)_���Jw��	}��i:�� �#���I�?՟�B����S�て�uNN�dk�R��=�Dq���|�<I�B���A4�R̺W�=�:�a���N�5N�<�wՂ*>�@v�zP����$����J�a���V��n&��iL={},慼XXZ���a}*�_1k�o�/��"���M���_4��KQ=G��墐>^��H��+�@:������bnH=nU�����s�Ώm���͢�=+���pv�Bds�Fe����ix�E"aͧ����*@m�@H��,
��G&�t�27y�,����zݠL�T�-�k��w��$�s�s+����)�j;�u&��f��K�+�?���D:xMT�T4Ϥ�&dP)+�[Q�;�O�rG��Jx\��G?���f��6}�i��vj�<��5�A�r��9<d��_��Y��uɳ٘��`��]y
3,�����x�1H�d��Zx��
�|�pI��	�G?�)�6A�K�y	��.R*���?��Mk�x�Uq\)SőyMi��^���!�*3lv<~�41O�=�d�2U� ���T=���R�^+�@�ܞ����H�e�!M�%���4\����9\�"YȨ��E�6����J^��u/�ݼ&&;؟�f+��z���/ڀ�"	KwWr����VVY��e�G�� >~�4J�Ϗ�h&!��R��J�f�o8UP�ͦ���r�_�E��6�
J�
d�W�3H�l��J�Pߵ+���T);[��߰"yW/C��S5��CZ����z��t�X��p���\0�v}w��R K������61�$X �(Ńm�QB�	N��t;UP�Z~�eZ��(�B6b>b����eK�}��Y��#���k��su��T.u��UG-ݧ�O����I&�l�Zq8�p�'��#ۅ�gx����v_s�Wtzx2�m�0��.�jP�Q��X�� v�ۘ^�m;�HcϚ�yB�K�$1N��^*k>�����%�ZF;�1g7���1h��M!�9��/d��v�����`c-r9z¼������,�OI�E�蔦
��F�u���M�A�URO��7R8bʐy!ί�o��M�_��SJi�%�n9��'D�9�Y��R���\s�GK���*�oz�A�H��c�_������m40��c��I!n��1A��bD�kN���P,-7�Tє����
C��y޺�Ҫ���K5�p�\r�@�\>����^ӭ��1�����z2����9�$3�U�������
�~y$^Y�9�7gwQ�p�L��A�j�J��!���X86JU�{����o!�b-ӷ����� ��Sf��/��%�����t�!��.�T��#me��@=�8�^���=�X�O�]�����"�`���1/����R�M�=���|&���L�l�L)c�(�N��2�d���D_:���DyrEc���	x��\-�(��T8�dqh�!п!�pH�J��cI?������'H�&�@�$lm<�C:��0�S�M7՞5!����� +�l���*+���ݗ�m9����+ġ�_+��O������+ZX{����������dMu�˰h��j�b�;!�^iN%���"HdFI$�����0߷?j�d	N�:2oe����6����2м�x���p�j�:��Yu�~�1���ӰR&h�E �t�O�/�X>�/��zw��R7=����]l�9�k��z���)"��_4�w��"F���k᪤�8��{sZ&9yi���]���i�ɄکU��N��7���\��k�	��c��1Hwņ�̑�f����u�-�"�8K2˘t���4 ���'��t�0)qL�7b��}���[H��M>D��F�����:�7KV�(�Q5�����>��g�<|�8� '���;yj�qypL� �����d�}��&�W6�Z���/����߼��R�C�#|.������/��ץ3�V���-�6n�lx��7
���~=}#�B�q��r=E��/�%3x��< ���Tk�5!<M��&m�s���/�WYP�9��T���V>��jЄ(�P��pJm�����m�È�h�
Y�03�Q���k �I%��-�G�E����^��0��DTyAL7��s�OL�	�g�h	��lz�`�E���CX'�I#�4j�L�3�k���k�i�q�\�$�M�G��>}�m#��W��zOҶÁ�Ukp.p�8.�G`X��u�[����Zzl�J�^i����V�8�j2D�9�t�Xkȴg�n��ᾩh�s-$v��E{'zs��m3�.����gY]�φ!�܀��/,0k�j3z��_�(��Cm�ᩕ.a��'��p��%�=%���&�n��{������Io\Z5�\��+��b�L�܀p����r�d�"O���L��'�+?��^*�A�U蛼=.�8:��T�8B� �s�(2jv� e��4�������B��cpd6|�X{H�^�:�__�j����9����q)r��V�EaJ�ܶ0+o����<o�˵�9C�����j�e��2��h7$ܵwō;�B�Q[�F ����Q4�>ъ�"%?���Q��FBG�U�aw�q��g�Ͽe;�U���c�6P+26(
B�ai�}p��K'Z��%���Şy�^A�E�~`�`�1�!��n!������'{�}W�gڋ(�m�y�\Y���T[T�;�O�s���\�Qz�L�$8/ꎉ�(��f�o߱����.���i��!�����lx]W�cO^#�I:����0�@������=���v�N��8�����=7u7�t%�EA����4wh�(X�ɓOU�x#�$:@���`.5(��E,���E�-��4�/D��뗔1���D�[���V��V��_Rl�7+
�J�_d��a ��^<u"��*\�Ĥ� 1bYS���C��!�G�zq%Gx�j��V�H|�������,Z�Z7�a$?oP$�	�JU�W�e��7�oܿ:6'�$ؒ�2��b�! �������c6&�܊%��$arD�BH0�v G�/�əPV��n�pX_��;�=0�N�(~r�I*�Q@��~��F�@OC�c"'�	fw���r��'>H�j�F��C�%��7^診�`ZS��j�0����"4nA�.3hE�:���Y��� )Ehw{�V�	E�Y���^S���a7�����R˰�D�m^�~�&��c���a��\�J`���@������+\�u^�m~�4�.@�����X�@˯�.d/�ɶ���<dZh��F�y�
#"�Q��X���P��?�}�#~WUۃ|�>�89�Ħ`vi�3�"x��&�G�.nzmM�aYv!#M�J,��!>��3�e�@2kGge�M(��l5����[�-��^j�!b����!T��tH�]�I���Lg�g~1y��h,�VQ.D���M��e�&� ���^3"��E��֨��)ߔ��y��>܀�Y�� �9�T������9�߂v����Eqm�WJ\_���	���l!�W G0M�F�_+�Ͻ|&�E��]���;��_@m�2c���g�5X�`�+�av�9h�5ؖ�"qm&oJ���SN�$z��f���Ҧ3
3Xe7�9������?��3� �a�$X��frrX]����mWf�7�W��]n� �:�Z���6[mФ���\��� �"˰�`,�M�/���3%����zŲ+��=��R_��k��Ly��A[�(N]Y��(���g6�T����]��)�D��_Q�h���L�G�7o^C�?��i�p�u����Y��{�,�i�r�L�:�[i��	p�sD�ɢ�Nc�������ܣ�)�S:V�?X[���^�ҩ��=%LǑ���N���ڭʟjV��=B�K�Nmc��w���ԊԂ�r;�a���o��r����i8�����"溱�E�:M�#<�HcVﾁ-���I��!.��$�9���9ߊ���y��I�&,�G��s�f�*��}�X��n�&L��x�H�54����+u%�y^�M�;��[���C0#:K_4��{�)&�dg���������5�lDʝS�o�q�.&���w�IG�3豜����/���=0+�R���=�Ce�����f�ִ�%ў27�}r�Uq`���)�#�c�����lw�_{��39��j~��8"1���K�;�5P�҇e~�HxA�%YV�8�vc}G.ְc�J�:��ə�izo��!<CD���*�+��G�O�xv�� �"+��E��/8M5M:b��ɘ����達��~;�po�m�ܒ�қ*E~���!
�u��!1̥x���p �b��l�nH���mVk:v@�t2)��j�?��ph����G7�fr�#K���l� 	����y�6g׭���'�b�Hc1A�_13K�Q�%�P.�75}[�v�a�\�����	Ү�x��T�x�8��)�IqR��&��h��������4�dӅփ��}��@���R2��SVoR�#o���kv���xE�HM+.L���dz�r|�v
:��!�"D���8n�ֹa�y��:��y��<����L�y��-���-��HQ:_s'ݭ@b`��� J�?�������|3�C-�:�"@	�� Z�c����#�]��I-�4��;��֎C�GV�c�J�.�95=�^'R8�v�}T��SW�*;�
m�6A�}�_F�;JTi��"%A�;�(��6��:��bh�+��fJ���E����y'^S���1I�Q��U��-3I�,�R�T���-+ڣo�?`a�V�B���k�z[ ��n?57���ͥ��ȇ�8��Y��+M�M�If��i�/����X������֡���]�<��Z��V��"���r#>�/�.�d���1�c����N��C%�C0)�1:g}{�NA�������&S��l��Ҡk�k=���z�Ų��Hn�&Q�c�R�����4���j����銩�{T�wI8���/�qMJd4L�y'�Z�Q��f��	@{`Q�_"��'�/q�T])�|�$�R6����"��B��&����@�j~}Ω��ߠrY�uqU�g�E1���n�*p&���K�) l}>���>���/��8I�Q&�/5�D0��i&]rku�������s"��؊l�Lь���_`h�T~|{F�{���<J�p"(����䤁@t��Kd����#i�G�y|O�V�Ʒ*�R_$X#������2��ҫB)����Z�Q���~��ۘZҟK-�V���X~�����'�/̰��=�D�[����~�`@>x�_�Wv�W#�(h'�]�{�a:�&_�EI:����7��<����1Q��ײ^{�܍���VW�XA�7��f	������oVS%_1Ǒ�s/����cG=��IK�g������a>H�L�|RH�@ �U����֪e��.�f������z�_��B�{⻄�"}�
s��U���X�U��]Ŵ���;]�bvĦ'
Eh�F,\��j��ݲg�ˑ4裙�L_3�U�1-o3�B��t�g�y����n%�847���6Q�ȈV�#WȆef�[X�n�x�T&;��z�s��ؓ��ff^��w����BI:��&��Z�j��'�;z���;�aG��Q-����6ؤyz�e�ni�-�cwMl5٤���uK
U)Bs;Q��Y��r�/"�=����善���/�H�@6^8*(��)�:���X��.W����y��Y����fA�[��c��m"@^���"W,���	b��-9�����Kx��A��S���*3��B�7Ԑى�O��/Nx�Δ���+FE�|�r���!K��\|�C����c�a����B5q}�n�����M���",��_0� � �VB���B�
�[���露{���??��ֱ��w�6�X���P+T��6~+E3	������ԩ����W��]���q�-ۦ͓��]���C�C��D*1c�7�ؠ*�д9:t�w@�q,[.��C��`�Gc���%t�p)
״5�d�����Vlh�J�R���_�8�΄Wbo6��P�Z��A������I�x�h������~Q�P�ȦK@���O�*����y1A_�B��j���H㶞'L|G���COI�HFu�T-2%_��.'�x�
���N�.`��]���Cb�j�@�W�ᕥ�V�_C3_��}W�1�,ǠC`�.����k�

�׆�4�εh�����&�O�q�,�	������ĝ�b�9�v�:��R�2'X���om�v};��h�Jx�0��R�@|����Q�D��0�@��Œ��ad�i����ͯ4-�M3jU,-�׵#�/�\�����9SZ��Ps�V�{>�u���������2�5\m�&}|���ֈ������J���u64ff;?�ײ��B�l�L�B�$�s�u��"�>Q�_Ʒ[=�%���P$_P�Հ)?ȶ �u�~�b�`�:=�_<���O��.�ݪS�?�+H�VH���@�Q�?����<G9.����d�s�x� ��	�QX�G�9?4��ƒ6I�;��]+x�gn���f���;`6�ԡ����%n��J �#�W��������abh�o��#9u��5O
���gZ0��-)6�y�姑�=�)��}^���J��"G��p�[j�*�w7`�+���E0���h�cX-0�͔�-1B�|ag�Y�v鼑��:��iS��f��B�����������3����bZ�r_�#�s �3zB4��QӛH�J͹+K/HFӼ"M�2��`{�_�� ���xm}E�D̉qb�ˀ�@zjS�8���JW��B��O��]��s=UP=����UX�NT^]{�.��Yζԙ�i��|�zrz��Fz�<F �z�ML�c�i����`�_Y{���yꬩ���A9q~��;�4/�~��z>�}$x��)�S��"�6�������`��� K�X���z6��CbW��҄$�>t�D�vU3H��(�_ds�9�r;���p��
�S��)�!6��A8��1h�qk�w��<ɞ�+Q�f�X�L�m���Jz�& K$#S����˼�_)�v���~S����=�c �|���Q�1k���Z�g��S������"��˻���b�>[/=jݢ�L)�E��Mn�t��}�血�^��V�S:� &J�Z:�Q����ǎ����
~;�%n2��F����{��Ƀ���V�:.<�J//GP�� �z���-��AFqh�*�cV���Ӧ��ӢehK#@��n��wĔlH�r{��$ƛ��W2��d��'M).�����"�@�{t�~�J�<i� �Ҝ�ޞ�xvc��}:<Z��+�	
&ֳe�7��:cL�H�����p�#��\6	���5�O�P1Y�[�5���.Kw�ϼ�%I��R�O�e�]p/Ǚ]_���(5~H�,�<}���KA_IC�G�ܓo�[��άF�DP#yr�T"T����c� ����	�UIl�J�wz�y�Ѭ�,�V�Q]�1���W�2�8�
?aX˄ߑ/��v[� ��ǍJ���:�c��(O���;?_-��3���//w�Q��@�5QmŸP��+v�ڐ���������t��P�F�'Cjb�a�{A�.�����L���J��H�&��bS4��9S���c����Sx3|��H�8:����1�'b����~��l>��Q<=�����ke��v�8
��]�	�J�g!k�fl�o�Nč���cfG�����
QK钑�n�Ѱ���G-|Q�1�����S�Y�v�����|W����ej��9w-����{3��>�NZ.��m;`8�̇ꏟ�Vg�=ޭ�@�<CR�X� h��R���T�ɫ>�����k;�̎�N�t�V���W�0{Bo���!Ւ7�F`:y��W)�L�[��₭XI����������(����zU����l�E�c��~@�_��!y"a��O�p�X�z���.��p�lI�/
�g�-aA~9C��,{����kE�S׮��a\5_9�;�.�g ���g������b�-���.X�좽��"��.o�ߴ��m��_�W��cfQ~�*��"}�p���H�'2�r�tX��2bB���N����&(��hl(���)C���"�kN�[{,�����0 9)^�}m�$!\E����!ǿ�r��Of�5o�6�O�^��7{-��5�n�L>�$�Y$2�˹���!O�(|mV!��0�c+ 1�d��B�P@9�J �8�ٌ4����ł��.��8I;	��N$��!��߮�Qk������[�;�n�m�w���C�1�0��lM��?��T?)�>�G�g�Zؔ�<K���X��^��l-��r1�)x����F����_X��B�V:Q�`��9�-h��RG�������6&Ǧޙ�ͥز/�:��S�T��C`v����o8��2�E`�����v�������y('���B�0����ٯ{��&ppV>Wv����� +���>N�S�%?Jq���apI(b�;��샥ɥf��H���w�4B��R�&���zƜ���3�ȅ�,�n�;�S� L#��[�\G�C�a�p�e+,��)�֜��=W9L)$e)-�^�.H����|�i��f9'�>xJZ#�A�A�_:�'��p��?Q�v�����WX䖾�3��h�bB�c�<-ل�-�s:�v�_�o�Ѯ�G:�&9�d\a鼔�%}�ɋڰm�s|�Ԕ����p �4z��}�u�e��@�ɡ��ώ��rxPM�����	 �;Jց�-E�o5�[��,�W���2/�)����ji�V���~:���s��=3����Ӡ��ks5rn义��"����(x��f����yc]���Jp" �H!Jնi�R�KT�ć!�?1U����=s<+pU�-u��T�ۦ��d!Yc��}n�T#��A�X���G�\�������®���S;�#�I���2�lX�O_Q�Σ�=�(aV�Tk�Mq�}�`���r9ǌ��X���]�'Bzg���NHm&��uH�bnG$�͊T�[���
#SA�⨍��7i�tN�X�����vH�@հp�5����&G?Q骞�(��*�H�ҿ�j&E���>B,�X{)Hb��D�)��˃!_��gX`��=l�bz�e����ᢣ�~��oZ�|�G7~G):S��K7S�	V�V�ׯ�*uP)ʽP����("�?�v��l���Ⱥ�q�w�HpHr��jLc�Yf����ؔ���f�(ʅ�V>� Y�[����8[RcVh�¦!�+G��P�}�γ�
�'��u���U���0�w�k�pi�	~S��y��Fj@I M���/�=�}����#.�dm�=�p��nU��:5�bl���:�8����?u�t�)���P'��=�>�W�=�/���?1���kwJ����g<�|��1�ŜȸN|Ś��0������K��D:ƭ�-�p񋩃a܎���Ǎ�t��Zrm�Q��Z���AJ$��#�.����DāaE�h%,Y&E��q*�����_���Ҿcؓ��LJ��a�x�#���G��Ƴ+-r��b�g�W�)˦�50��3☯�ͰŮn������4jz]u�x�}\�>W���Ě��߉m�� ƚ7	���E�+�A���&�dH���Rã��a\ź'c����^���G�d�0����2����Z���Кf���r���p�m5��9�Ե���XE�i��G�6�[�;֊_D0C{��FUe&�y,h�.ro�i�ʖKH���p����Ri*Z��x��|��V�X�gi.�aD�"���,��&7�K_��Y�zB��K�i��Ӂ�Rڡ�[���g	&����/:FNOqXt���\������n��ˈ�簗�W`�(�?+���)�R�l�s���f��1\��Z�{Z�IF[1ܶ$�|fk��!�O	nHj3?��)�?�ݛ�����-ؑ����<�_ %|����,���rK���=�cT�̱����Lp�]'�,'����t�A���K���n���fv���&�n1���_n=K�j(�3Z���ᙝ+K���5c���j��4�������H�����Pu�>@��N;˄��g�F.�ăL����QO� ��)�T� ��^I���ŒcM�1��2$�{j	~��R�㻙.�S��L��s�X�D)45�B�|ꑅW�|��Ǝ���q^��1կ���D��Z�	�=�LI��v����d�-�ݶc�`~����)��d�oP��o$L�Kի.��'[j����u�丞��43���6���%L4���[���qQ��w��f�*.>8s�X@����? ����!�L�g�����VH������/3�q�x�Pő3�M�Xʊ/���C��N�63��4�m.˘) �w�K5?+?
� �qH�Z�bWl�I��f���'�[�u���	�Vޘ���|8i>��;(�㌨{ �����U��6���j��7���3?�gd._�\����* A�,fգ���X>�޶�Xd&4/�o��r�,���/(v+Sm<�.�S���(�߻�3C^�5�=n@�o @F�8婥8
��a��d��`����j'��y$y��,��[ �� fJ�$0s%M��)��4��X�=�m(�S^����c��Fo�/�5V�w��m�M���߼E�?�	ibl=�ޝIK������	a� _�G��� 3n%7������U��da�Z��8u9@K���D�"p!w*bu����l��u���/p����L�h��3���V]�Il�\��7F�5�1a;�i1S�,�:q�Q�U�xs1� �S<���1l�u:���[�*{�z��㬤�L����-��C<��A���"�����c�"������Va�M�v�UT�4�9�ȫ���QӋY�o�%��X}��3\�B�N+SO�A�#^H���W�C���~�߈I���u�W뵞>/� �KK���%���5��:��`3���3]�7�z���Ǡx��M���[,D+ɌWP-�/y޻St���6��Z
`����w+���Y�kZ+�V���/1�c��g��<BRϟl_b�����-�=D&b�<t���d8
��2��,��@>��P����:��Z�?^����t�6yZ+��t�:���O����*u\�jUΎ<�\0�l�6
ic0�5��2����ք_��j�{xb5̩��3�I�CgV=�ݷ��Sg��&���Qh�Mp3�z��Yr�l����-���]��N�)��V*���I��g������~֒ݘ��̛������y�/^d산�+E��q�\�YҫU#ǈ��J;�&��,�e�a[AL6�~sh�K͟�dO�A��pUWBBvC��S2�95�8�طp箒��Y�����	G�c��Z��p�⾊Z�,���Vs�^B��C5�!Y9(�M�O����k�dX7��-��T&d�R�+�݂� ;�'mI�X��e��W�t���J2
�U�S��9o1���T]��2S�QL�ko���3N��lwA��9BLS���Du�+�@���޶"��D&�4�� L���Q��v�cw�("#	ňP��j	�8���� ���� ���JD��^^:�jK53Lr7E�Z���Y��kCt3x�(��G ���`m�Ջ�I�Ac
܉���IK����On�d���(X����vRH]�����aE�|r�S���[�+��CH`�'��)���t`�s��Q�ڭ���]�L)��!0���3P����f���{���5>q�*~���\��#;.ًݖ��,���/ˡ��c�'�QZ) ���lF}up'}��v|NC�F�Y��-8�W_��[Pp���]����M��M$�	G�`$�7v�6��7D� !>�Lgw\Ȍ�!�9�����u 	v����@Pq)J'�������gl(�J�ZD�K����7�����#��KK�����J�X����ØqN���ÇїA�$���gs3�o @?zy�
�B�m��7̏�_��԰��(0��CG�P��O�%�BE�7�?VL	��J^=���[<f<[��2�޾�In~��co�npyA��Ӧ^>�&��~v$T%ݼQ�H�T39�Vؚ��.M�W�O���#n���wH1���Q_XeH�K$��7�f"�Fr����-+�?+�{�^��Շ�������=dХHU7�\����ӷ��<��d;�R���w��Rq$_]N�f��Ê�T�py��2��H�Mb�f"�,X�u��6Gl�@zG�G,.�3*�H1ߙ9�A��������LDx"��C��wUvǷ]���,�A���A2�,f�w4�Ș&JL\�<}<�cus����yɖz�s��ޒ�� ���̊$o$P+�a��tI�ε��hC�r]�F�Fe��_�]���{�#پ�AA��lkRM���xm;��˅��K0�����ˋF�4��R?�a��>� g͇���z�E��f�'fY9��T��'��uu'��yldw�g�	��T��b�ȟ.��=
�,����>^$սƻ8�sXGZ�YH����?��RMP��;�1/5���熕�T��k�䰗�"