��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�/Fw��x��b ayk��]���
t����jw-V��k�d<a�f��xx�/�~���)ҁ�چP�^4�#�Hy��9�=���
}na����ʟg��������lE�R�6By��������"'Zw����k��=y��9XmLjp�՘`/��z5 ��r8���˂}���\c���ô5�����ts�r{�ش�x�W�ʹ#[�F���\hU��5���.f���Sej	��`A2���r�2ss���$��޷VT��O�P��'�=K5���)~z<����]�N���9���<�����+�<��~�eVc��rE<�=������6�ζ�l�d�%�8zϬ5�T�ɦ�ڹ����Q�<�ՙ+$��ѐw�ݜC���͚����d>"�i(�a�D��ʈ�<���Y(���0���]u�Bh�'��Y%90����Ŷ�S�A�D��9��V�mX��,d�ч2Gd&��6Ba$(����������xÆ�a@a�f�_s�'�9�_�d�-ғD �)�1=�Ue~b2#��LQ��S^�f�ݰ�z�B�/9Q%6CO����@��nd��~�~Jc<�_�ff���~n�r�S���W����#K�C���Uys��tu[0W�@�=cq��2�w\�O��,��x�>�e`����T���ki�U�vH�a�/N!I��#�6�nKȭc�����n/0wz�"�r��Ī[d�i�zw)���#h�U?29��.�HbctU����jI�N=�.�W�����c�l)��Km�A�U�bhɽf�jm�|�t=�9����FC%�5�Io�>:�9r���U_�[(>�g�z|�����o�#�VlOf�[�����.�`f8�ۈ/�|z�q��
���mSo�%ㄝ�G��,|��9��1�����R�A�%y+A.i�򤗣�;��XrC]?����؎�n.��\_����*6�?�G9ʮY>�<D~s�j��������J���4|`k�ӸRCDD�k��,��K�fS��2f�Et���R\l(���Y
�
��.�9����*�S@����ã�ǩabP�Ϩ�"�&�k��p��� z4��]l��)$��=I����������`.w���K-'Ԗ	�F ��c�ٜ �<IJ�(\�#��v�4�U������¦d�6�l	.B(~�
�Zs�W8m���TdT���H�%)'B��O;�5k�s�:�����%��t�e��F;��^�Q3�v��4)��t|uS������ Ď������U&S�̼��a�z���O�u��L�o5����m#���}N�g�u4-4=���-�0�Bڧ���+8c��FUO���I*�Z�o����RZ��;2�,Ζ{��WK �E~BT��䭁[P�ݳ��p�R~̦ ��볟��������־���^� �()|��4k
���RXQ�(~Y����7s���3�ݺ[�<�+�0���9�B��Z�	Zvp��sI��.f�E�ǥt�0�W�.`� P �A��J�/��Bb��
_?d���'gr.�Rs���dd7̑��R��d�zbz��"]ֆ��������hxr��g�f��ʒ�K}p	炭��n�6EG��:�0��*Ϛ������Rj5%a	�0�q���}�'j.(4�_�L��R��-�(=��l�A�e]�M�%�$��ė����'�/Q'���$Ic�Z�`�b����x�d0�Pf��xA.��b=�F8Řdyi8���N�S�:�����E|��/�8�L���yʆy�3�A%'{H��h�p�/�����k�0�0��,4r�'J�]:�ƃs�W:4����n/���M��<�%�t�E�M\,����^�g�r�������Df�(O�u݊�	2i���LH� ����F^`�*{�e�C$���9��B�R���O~5�����n���^U ����^�K}���be<�D�F=_���:>Ai�)<�>�(mHDȀ�F@݆�����N���w+$K��l�(kW����)~�.ōk/�����j�/������; ��|��Ll����񽰶�"��[�ɴH2p�����<�`�M�V~-�[�3y=0n;%^k�= F�h�3��ؤ8�A�ϛ%�f��b�������J����)�ŸM���� ^����\����K�=��ZmR�������2R>�7\��ͧ��u*��m����	t Tx7"}���IbR<�֞�\��?�O�#�����Mrp+�zM� �C6l�bGa����K@Zt#N�[�7��<�[�)�5��I0MR��qdJ�<�^�HOx��q��toQ��WŠM�w�jh�mr�����o���t m�������;��?�u̮��|�L�۴gpW���%��ϱ�-v�g
�-��fZ*�F��mƱ�>����g�D*蚶j��X36I<�Z.�p��W9�.S&9\���$iR��(=~Xh�8C+?���+r��W��+:�p�#�(�
�}aJ8I�O�C+�G�l"�����2c|�nF����6J��/��Q��<&��� ��O(z�A{N?�߳�P"���6���ǁ@�����$�Ĉ�%��xr��TX$�� �eR����\�%��`nK�t����2%��ju��5h�]8�ô&c*Q	�}�\�WpW^G��ȁ����A�5�7�j:�s ��ס�:l�%É�	��{�5�4ܦ�y����^�Ba�ӏ�0�y=�����0�]�yi�����