��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����d���o	�i�Y��ǢNFKR�r�d�Pє@I��a�ڒQ�6�: �m��H/S�ߥ��x5F�
��,�
v� ���U�͗A�^��!����f�f�Lx����6�|�G��ӗ���.y�o�Ke�_6p�ʆt"{�oe��!;w㼒K�C���w/Hb�]�Ks��a6������`�P�M��0B���@�������o��:���T�#п��mn���-�6��9��3���qu�Dv݂5��q#Ѣ�.��%�}3/��5��#W�$�۩J�S����X��(�&1�nr��xǏs�'����{�&hb��P��1B��]O,�~AY�������j �Eۨ	m��C N��A�1���(�Ѕ]��d'P��v��e��to���dt'�9SXh���"m���_�cA�jj����d�+z�m�>#���[����Q���LIA�/h~��jd�7ov�Z��;��Fm�����~��|�3��*O`�,{g~�d�BB-�g[4�DW$�x��yp��[�vw�E�('�>��������jl���.��Au�4�$�:��m9E���ܤ�� �-�E�	��̶����l\K�t�4^�Z�g춿ŏ��M7`�
��h9j�GJq���U�<O8R������D)/90��vc��&P�⇚��c�w:���b����;It��:b�Guc��b��myBT�ޗ+8�V9�}+��rK�6�H!�B t?�����Y�E�B��m���H��=�ɗ�,��ի�c0F���F���]{�\�S}|�K��Y�����-��g����S�#r�=�keiW9��j���f��A���uL���>�Ɩ����+�ݒ7X�Aښ����$�����q��~-ft�ϑW��ԟ�l���6�7��h�e���C?�����Ϲ������Do�!���f�������@.N�W<'�P+B�E�]%�C�Pc��~C�񲟄V��^Th�Zm'����zt����N���Ґ���t����Ƅx>֋���ft��+>(�&<9l\8����5%V�26���s8!5�(�v�aF7YW�{�5����k4�ށ��Vթ0�DVI�pR�-�s��?�P�λ'ȃ�(v �_���D���u�R��ty���[��=VƦFf�w�"��VBqb���/3/cu�S�'bf/��O����y�5�b��L+��z�$��)�x������<@�[�eܔ�ERA�j���V�5Ѫ�����H�=�����r<.W�X���V�ܻk]�0l���%��9��G�G�m0��E�V2P~�NͶ�d�,..U瘅��JZ��Ϊ�ټ<�.McG@,c/S��1��݅��mlP>��G���~��b�vsF7��ڕ�9����v�$8O@���Pr�Լ���9���A2�ܷ������&�:��(gv0���I��czϚe�H����-��[q�$ �E���<s�^u�xM;��cӍ<�!�~F�E:�:��0��?\$��W5M�>[�wc1�DV��ah�����9+/�\��7���9L�`mm�.����X�͇�+�Ŧ�4���;s�+9�V��O�F��5�W�x<�@�$'7U���|��h�F]|h9���(�4��3�J�+֒���YL�h�����sEa����p(k%
=��l��ߊo �r.�ۦf���z�6�x��Pn��k��������[���x�ͼ�0�L+�Hc8�(b��?l��|@�"�P�%)� ���Y�>K��_����������_�8�o�7&�io~;R���$���l�:
-/�L�wpx4�4�-����F����N6���)����2n�c,E7�O���A�&n�G����ظ�ئ(L�R�,��|o��^�f���-�(�JGy�Ei�g�A�0� t�zJ�U@Y���8�J�Y�(4;�zV&	�%��QZ����hs�T�J�P?�Y�D���>�03�nc����Q��D&�����ٯ�cs����
򁢻���c;s=��e�W�T%����,��k2P��Pm�"p�f�T U�	�xо�'���N�t_-��|R�;+3	�*��5�S�}+���������!���R0��EAdGYYS���#��4e��������<"QLN@���v��
2o����X,�����fϨU�?�T�(��b����������[=���/���eȨ���Y\'��ĺ��&����D�nD�+	N�	".U�YJאt=s�ˋ���Rq�8Z�dMG���NϷ���$��6\�Ky��)w�p��-��]]1�'�E��g�-܃������z�X���4S��-����E��Ʊ�|��?<'��J�JU�?'	�B.8\�� �ԃ]8X�>B���Z�ZWG�YRK�d���vX�]���J����A�f�X\������R&��,|U�u�+'�V�ş�Q/m��f=�{TZd��}�_����r�UA�&�cJ����X�1n��w�<�L���ڦ-Uo��P�"Iո��/�w5kⰓ;Z$���	#�$<�7|��)�P���zM������뇅�w��
P'dֱ�.��Rg��" OGXV������Ǳ�9�h�yŤ������ו\��v��Z�%�5�㼤E���ѵޗ$��j*�b6$L��NU�嗮V ���97� t�¡ú�8�,�1�^�2���m��J�E�t����"=J�g���sNq �/���#Zl�ho�S��Ϫ ��,5P�C�{�Q�N��g�]�Ԣ$A=�����a&�6[8��j`,�� �o�Ҡn b��'��iMR���.8�^�Ij
	��R�v$�Ƀ���X,�����P��J�h�j�ԥ
B���;�c��}Y���0Ŋ�mA�s��a�k��9�F~r�˪��K\Q�߱�%�(�����2�ʼ�Hs�L!+.���Wj-5t-������2I�Zb���N���L?�K�M۷�"�&@\�rg?	�Į�˓�͟1��+�@G�?�2�l#MMun�+��=9��	$q�qo�b@½(���m#5IR$D�#I��-F���J�� � R������}؞gm��^&d��E��m��F���,	�=������p�&�vFbg�Ȅ��4�]��e*�Y�.�GM�B��G[l��֐�j�-˶�-�0`�])�����*;�\Uk�gP�[4��#�u����t8�Z�E�lwSd	��r�ԕ=��_0h����E�S����)�.�K��!�K(d�v�t��@coZz�Ic�W��ɿ7k1��ve|�m�A���qp5_T�o���=e`	���?S��o�b4�@gM\iC=���3�1�"�'��w��`lv�
��A�%>�����o�zs���+�m��=̞1F&�.�v0x6IY��~��V�H6O�2��Ѓ�pJ��K��jώ�K�㱐�m[��g�w�q=��̕˪����q���IwK_ܯQ-��_��툥��{�֖δ�/O[����h�leV���x���x�ec�1���& a`�&*+�S*�E�P����Y�$N��|Z��FڅE���>:���`����Y�-���v�k[0��yg��|Y�?���-�-�c(���0X��xG�g:���2D�rX������w<��5�($�J����Ų��d'{}�|W^��ar��7r�**X��DV�)���X��[�K�C�	��e�A��ņ^u=�F1�Kʘϳ��.30ɫn���}pJ��I�w&XsdŊ"�}t!]�W2�|�L�;v�%�*I�s�7��e�a�G�h:֪���&�����7��/�W�:
G�u�ϳ��m��\�0+�b���LK�RИ�΀{X^x�vH.�R�w۩X�f���c�b�
�����έ|�b�X��3��'e�$�'�B���Z��+;v,|�"\gK���-���aZұ���⭫�.�ڔ�� �T�0�)"�Z,����9y!�M���O�Y`3#�s�q��r�ZI���2�n"!Ha�5����&���*C����ǡ�A���Q��}{똢�wU;� �Ƣ�%kw?����KM�����������1m1��P�t���Q��70]9M��S�b�<���Mo��[)	EM��v�g��H4D�_v/�y8�����g�6�˼�3�(�C�ʝf��&��~��(��~�2�������-s�G�Na����HhMA��Ķ��^J�J��n���'��α}���8���=�o�݊����5�����^�a&����!L�ք��.�I��Kk"�p�Rc�U�骻�po�=�ex!�"���g>վ�̂��3���b�Lk϶�n��Q˔�M�ߣr�(ZE>��][�bZ�+�)S��N.��c[q�C�zkS��#�X�V�S�����g�fp�?�����_�q�k[mT�4)#)�oŷ��j�\>H��6�������΁8��O�5?ta�1��|{*i�|C �Y�� _~;��jH�<P��2)�8�Zo�L?��E��*���O�WP[r���UV�s�&h"��؄����tʲX�Rg��7�{qv�p����)�����U��I�^�_h��V��������Y���u>�C�u�9� }�g��]Md;Х�Bv�����:��P�ͅՀ>J�~{��f�RT)lfuH^*֨rW(���z�v��1���Ų��mڛ���0̸��[Y��S�������;�E큃� �Q��`���4>G�4x[����h43�-��y0���7s�}O?��%I��j��@���n�����W���w�A6p�l�xjtgI%5b40C�g\����d�Q)jH&�d1�xP��,UbiV����NnO�Z����6󐫉"X�oa�� �H2H��0p�p9��_m��*�$�_�S�����va�O��]�n�"K�G8���'i��*2�)��7,ǀғ�!��{�A'�r��a�q��exT�z�$�����{�Q�i>^%��g�P�F[(00��L�_7y 3��b>c�Ҩ���]�74u��YRȅi�u�#+����2��g�`E
0����b�Ud\<��f���9h=m��C�T����t�}.c���E��
�P��^1 ���{�����C'�����ʋ��=��ĒGx���w��׺�賵�-[�c�o��<@ģu�׏��c������G�[��'B������b@Q����Ȏ��������(��q ���70�jiv4{)5��8��v�^�G j���$~��rto�m;�M|�l���O�3��:�ol�����;�X�����皵�]�&n�\G`~>�QjA�v���QLD1�K���ܑ�{�|��r,K���O�;}�O �p�6��W������r��Vr$/ꂈ�W�uF|�Z	��b�F�،�G�:���3�<\�=08��nQ33�HӸ%��;��y{���,�Mط&	�3>�v����������J\������,&��w7nQ��6tR�!��'p�����j���{��P�v�	Z�;���]칁����}Ԅ@���pRQ,��[/G"��[N����bxˢ����z �O��5�jێl~R:ˡ#nr��,ĺK ��V�0t(��-UH��-���[�|B˕��v�8�ʗ��`!+T�:����NoA�:���l�ֳ9\v��C���d<���l�܉/���4�컾p�ܒ]�`�7|�+�����Z�"!�� 0���b���ԬW}����u�с6y��ܭ$l����d,Ǚ�#�Ka(`<0k������8v`�5J�f8�7H��]Cl�xےߑ�nRG3���h��n���� ڕ�~��v�?u�)!?�ˏQF&���<I~�5<m2 �����u�r:ӃN=wC����Ơ=O{	z@�Ah�Է��x������=�&'<���U�D��܉lhd���ݶ'���!�J ә��T7{��Gu�%̂*����L��*~\���>�n��H�Y���{@U�p�/����րm�x�\��x�Z��6���A��(��a�VF��9&���Hm[�fC�|q�B�9o}(��BC��k���X�?Š�g� �J4�4�'��J�<>�;�t�$�UW}�F9ت��Y5�K��ȵ��y�:�B���ӴS�Ώ�x+J4��Q�V��D9UrJ��pP �h~	Gy���<��w��uS�F�����\h�TV]�,�nWOJ���y��� 0�Z՘���].�;�b2�I�M��3(��۵�F��]���``q��6�B��*��
z+0�f�/%��<�b��1�^�����
�	�[���e�	BL�7^�������U��a�Xʶ��+��d;�-�\���a��ң����4�^�P8"w����Y=��/�R���M�i<i�9�N�$"E�^��k�� ���)���j� ���g9YC����	]"������eX=4��ɝo-�4�sۓ�n���7�I��;k��4�녌��|"e+�@;-O)'��C^�j����tE�6AQ�gD�3+�lz!���q2�8��:�y��Ȟ~j���%�2�S� �)�%/��bDTg�j��/���=�tq�]�7�FYINɡb�/�O���5�2�%1:�&h�#�U�J!��ɐ`��p��
YѢ���6��k~��a̛�A���T h	l}�T�'���M哗�e�礈U� ��V� �U�� �5���9\y�[��b}�㩌ۃ�TIQ�[�����K�,gql�8�Z��I0WF��m����z�2��5�&��8Ѱ4�Ds'�"��B�Z��hE9l����Cr���-�=���r�%��F��m�������IZTC+�U>�2ϧW!��*1�"����� �Ό�3�6*jBl߅Qܱ�m��뛇ՎsQ�'b�S��8���Uَ���s
�d`�d) :@�N��M�+�Cq1�Pu��!JD�VaY���,�$ֿ��o�3N�bIU֢�x4�`R/b��JM�P�FJ��yҟ�<t�%n�8' ��y@�TD��dH�Fr�M�l��/��C��	��D�����Cj��Cǋ��5��؏�e ��I1<؝[R�,�.����H�� b#��lӬ�@�!�k�D4f��K�jq�*Nt���D �V��2Ҥ��vZI�H�G-��� :)�&eL��n�q0�y��{�GYR�,�Q���9n��7�TX��( V0x�Ό���
K���q��g�������KG6���L|<�5���? ��)���p����}��{|!(��R���ɿ�b|�p�6�o�+��?Fܨ�:FMZ��Ӕ6��dp�Y��wⲬ�AD
�g]J��n$H.�$P�d�`to���|�J|zD)�[��qy~�l-6�2�k碤�'�2���nˢZL��=�k�C�d���9�n.��R��ƫjV�Q���'ã�{���i%���əA��a$�{�� ;CB�ːf�� �K4j�6~!����"T� ������X#����{tM�i(���l�5K;v������=CIC�z�[G�l$���¯�t��xǑ�1KM[Z�.N3x��q~�g:�*��e:��܎�(�gۇ0��m�o׵�}��Ro h�y���Z%ɏ��
��6�3"֬e1ۙ���ԓa������ʨ���1��&t���@�j�הj�����G���$ܲ��k)AK��b�p��Ά�u�7� �;iVbr�[<cv�Ʒqc
��:�?�`�D>��s�c��و�;��`�����+,4y����^3ނ��|·4�t	̪���u�fG��/���?��>��)�6�����Y���H�zM?x��
�kg? G�{-��)g>N���V���wy���9b�Z��������@�B���e��֪O-H'�ǜ������r*^VBZ�������O8t-�p=ɏ�h�i�3�dL�8_Wh��ۛR���8��Fۼ��v�c%�ѩ�@�ߏgu��\d�8���?�;�������o�P�w��` I���~(�B*�ѱU��=�qa�/���Y��[$�I�U�ru�[L��w���.��M3v|����B��0�zn�c�)�w���G��T��'�;�߶��4��Rh���B�W	^�((@S�C�3aC�ebw������$.��!~]� `�d�!/�۸9U'���V�a�����Ò�P�X��)��\ER܇��$S���p-<^���]%력��F�2�:W��{&ۿ|0�>>�3ЈPS�d�!���̓�澃dKɄ��!}���#?mb ۱��Mu������ۇ�f�A<�I�������Tܹ!O�%2��᝻��~��>���)�/���T�"0�[fԧ����L"��06gG��0�b����x̻�2+���:��=��.�0���0B{�Ga�=�k��E��\}�Sl�����HR6R
�>2�@����(-AOh7'^�J#8�H=/mR��ψ7�jG�x��6d迺I�Q��L�����L�U������	j]e�5�p���$�H�b�QՒ���)P�M���ml���u뿨}X1�ac��'G�vYN�aK-�����i��5}�= ��z���u(�\��$���P��w^�e����>��j�se�������t���1r^��D�02-�H0,u�GK+\�7��8�f}� ���n:�ۀk���N��J��U\�L�;fl�%$� s���`/�����v�$íТ9I'qbY�!�\���~�BYJݸ���5�+�ii�@��]!�KIP;F9�m aoH>�Pq�.Ri�����@�T>q��/��b��/�{VUT�Y�"%˙�}M��kz�D&���3h��=׋����H��"�b��Ǵ&Ue%g��S��16�~4>H;����X�L�T�t��N$���Cִ:�i������:���إK�5!�4
1�n��4T����̩�J�ͳ�+�`I����4�l�S`�%GhH&m�X�u7��i9X�u�}���r��;�¢:\���(o�QAPH�t2�g���K�~$�|�N��b��ov
w1I�צV����kDa�Qv����8b��0�}��X!;)�u��9|?�h�5�t�H�z�ew���Z�?���[2nӺ��8(c ��:T!�g����T�v�񹁊��nJ�y��m��Iz� ߭�+�OQ��c�T0�J�I�n��Wv,E�������(瀮]�]�7 #g4�
�S�<��)A�e��N]��``��$�A�:� q��K�	Mg���|A���wG�x������< o�@"�^X��x��	;x<�@JA�Q���/��%���e���þV��>�s(�;~y\��{��a;+G
/�r��R���o
�����^t|BVuw��W-缐�����XT����+ܩ߫��i��g�P��uG	:���FtT�����A�r�QH�"\z�o����y��~��C��AlcS�e=�J4��}��ڲ�	�%1��%|����\�Xx�3I����YfX����s����X��f0q0�1k��!���.;ta}i��ڞ�u���Gfnc�>(�蓃�Ph뇷����or����.[����������q]��uw���4Y���xt>@�������q���[8�J��!��V6��Oj`���<��^^�N��Ďf�n�N��1j�����dA�E�� a�At�了Ǟ[�_��Bԫ�� ѪޓB��Ж&��pXĂ%���M�¬f#��F6%��Wx3ߧ��$�;~@��T{㕓y*���+_��|��>�cϏ�V��M-��J㯳򛕤qCr>Ҟ�O�/�����N*֡� I�t�C]�T&8�1�������$l�K�m}p� �ѐ����<��°�u��>>����V�A���)��-�|x{(���8K|ś�o�k�����ć�v�`�=vG�{���A{�l��l�&r�Ǻ�?t���[1��<i��)��Q-Yq�K�'[�ր�R�f�zN��B�� �/ %�۸��z���W8�yM
-Fo�q�M�m���P�90{�#
�h! � |�n1,��cMU^�t4O���4SL�nUQ9�I͎�p��1⬜�m�Jd�0��'p�V8�e�iQW9T(�9���;ʃ�%y����Ч,a�CIٔi���mD�'[�T�|�s�`�ps=f�]7�hL�ܥ�U3Y��T�2$�oc3~k�&>�Qt9��p�׌ixK�]��9o��5���!�ގ�u�+��^�\�+���r�=�$��h`�[�|�	R��{���[��-�V����
"?��s\l�AvE�����J|���
�����`ǣ�e����i��
;Ru����4��7���Ci�~����g�;.R��꺮��=dg�Y�Bp��8,z�P��|����̅tⓣ�K����Ju��V����z�8���7�����ԦCh��,�T	E�K�F�{m��(��w���KT�����}�Oz��'53���s����ːXj����=��+�刬��h|öM��y?��F��{�d�b�����Ѐ��]��Ś����ѕ������{B��%�0:��t"Bg����B�U��Z�}�ieaǾ����\�֡��A"�`졄{Oѳ�]<��-0��6]NsR���@����𣾽oJ���ݣ��Lu��W�e���0�<`�H�y9O�_�1��]�XAg]�K%��5����R��2>������lT$_�F:��.�f贺��J��G�&iv��`�������rg}�PჅ1x������eqH���n��s�f4��ړJ1s�]�`rE�<��Ct��WK�7`�7�P��v�1��Zt�TPvqg�lP��3p�Ja��\��
h��
B���,�#Y*m����]*C���B~jC��9>6+y)��>�ʊ[ty��z6�g�^�)���29�ǽ��I�n�坦�zQ�F@Z�cw?J��� ��*�FC��p��g�Q]]_��2���ewyE+�����ñ޺�Ӣ��51^_��!�)�ecX�2d�6���e�`7L^I��f.�DĳL��uX����l:gq��5��|%#��iұ�g�$�v�-M�P��r� ��;I����i��м@w���\��哪C��; ����bG�I�z,���7��O���������� �t��@�&4m�K�2�M�g��Q��������Aýl����~�i�'m��#^>�z	��5C��ȕ�N�N�k�_����'�+�2�:)�-�Bߡ�;��H䘌�,8����!���T�_�#٤qU`.�6�3iV!WhO���o��������t��z�:u1v��XM3�8�m�ط�$	(��o%�S����w�t:t�l
�������2|J��Y;֯d�	v}s�eE��Gm��t;�/�e�m��.gG���]����*�B1tb�b��^�Ytӫ�R���#�V�5��%��� tg[CL�<#��9�s R�(XI���B�k���#G�P�l+��Z=�2�8TxQ��7|0�oM�59O�P;\���?�ŧ�oU¸��u��S��B���!lF����Y���,~��>A+OP�h�lD]Z�IB����ځvd�v�����6a�bKd���Qo@����,;��¹��<x�j�|�]����I��Lr��ʃ��~�$.wD��êU��G�V�ҿ4�����f8��g�#�Z�CSӟ`�&o��R��Ʃ��y�����q���:Ŗ0D~����ߢ���K&Ig5e��D���Eu���g �O��� �����mJ�5&�|m���K�]�d�Ŵ_Z�g:r%v*W��.�/қ��^���6�e+9&��-ٳ�~��H�', ���Ņ.��	���a[��m�<�8'uN0�����3$��µX&r�'�>�N[��>���~�Ч�C���������Q���'��u����[���<����M4Z�L1��%�v��}�U��-��&�\�@S2v�]�;����T�Z��� 5Έ9�7cz�.�[Ƙ���6ZQ�l�"7�S?<��̫����|�kt���9�w��+��nv�!^�S$�#�t`+��o�/)�9Ȇ0%V+���e��)BpU	�0޵��J��#��(��~�ő&���`�7�xR������JcL�1��U�f#�N6e��5��̼��0�������j�l���r���v�ׇ#N���u᳒s�M5P��u�����0aݾ4��Y3K�F��V��AA�4�fJ���=̗�T���d�N�ѿ=�"���8{N�PC�:�a�rNK�|������ϊ�R�E�Ӷ	J;Zfp�2���-%�}kp�m��|i��Y+���O��H	»����%���ʭ�р���15� ��� �&��h&���`��k�b�{�eStZ��IW�F��)ǉ�
=	Nw��g�rZ�ӔJ����H&�����2�)���V�:�����?�ax�q��\�~dlع�f�4Osr����u����D��������Q��!S�S�]`j�9��Ï���0O��v۔�XA�8]�1gl#����J��"}��*���T6�䤪��]_[��MixLAffb]qY�"�S4.ȯE�;���WZ�1��-@��[!���'�{ �sR2pQ0o��B/=7�>��b��;��`)k������Yi�ab�%��C#�S�c����q��H�ud/�>��ćg��o�Y�,��#�=��z`�z��pZ�A|�Ҹd,YK��e����vB�Q/�W�E��"���?s�KH��V�ʝ?�n̤h/����K�o�%-ZB�(������?�\���M�e]�$��D�;��U�
���j?�z�A��Z?!A��H�A��^�*㩽-A]\�m��T���<���̋��*g���>�'g�V���R��V��i?�TX�N$H"1	����� |6���X����D�#Vis��s������O\m�b\u �/Nbb��@{��іܡ�h����r;�����0��3�,,��h��ez�/?#}j��ێ����ۛ�d�6D���N��Ԝ�T!��a�a@վOL穬��/����hdãW�q F%&t���#����戙V�2���M2Go �M7U���
��qz���U��\��c���\	�� ���}�=w.�M��!&������F6O��a������Q5"�߂�7�=�hT)B��"�y�X-]G9��ڒ��S]j��zh�Fq�I�vd�s�U����B�ٱ����v=E1ғ�Z���� uH�pڐB�Z���߳'f;0�Ïk�������X�i�� �����B ��=E��a�ۤ1��:8g��ٰ����f��1��N�{76��m�˞�F���yD`;b�A�i�, �w�g�`o�=6am��11~��S�ʩm6�s2�J͉x0תy`Jl0AO+��5����A��~Q�D7���GG���Y�b�z�0:p͈���3��4C�"��/j)�2P J��>2����w��dY���q���t�0Y���hbP�U9�_a���Z��!=òvǓ%��=�x����L���~֢S�3�U!�y\3<�
 *u�9,*}���~-��P'b"h8�D�������1����?׫N�jb�?����ci	n�1�j����J9p�Ǹ�;Ў��;��w'���e:�(�Ν<��4/#V%�XN��C�Z��-�6aj��c�Ń�+���r�9|�)kB�-�Ul���t�O'+SO�b���-dK����3߭�r���8�W������"O&�9�$"{=x����o�df���F���Z�����U(����Ì����G!��hgQ/&yS憢H�QsQNSp?�yI*6S	E;��@l,�@���BW��7�! ^I~��8�i�9t�Yf�l)-!����s+uZ��0�Hǃ��@���}�m4ZO!qX�4�رn���AC3P8,�1q�i"�w=vކ����뚦w��e��}B�^�J{p��(��� $�y�L�쨼�}g���"���X(�`�4�|tS���S�Zn���a-^�W�����P��n�[��(�u��$�戉��u���6��ɂд�����|�H�F��������;�t�+�I���i,C�_!A(pN0��[�U�)cVh��i���³��wnc{�4Z���qŭS6w�GuW���9`�2�/�(noH��H`�̚�H@�nrV����ǿ���k ��/-��	Λ��G��_��~�^ć��,�[�1WϏ���6jdK�C?yX����7Q־T_tá����y��˞�x���bq1>[��Iع�6#���u�,�,2g<&[?��� ��ຸ��ܿ=��{�}<��i������P��C�@ѐ7�Mꨴ��xStZd�*�A:^��W֝�>�	�MϠ�g �4�C��S����C��s[��d<<E%&�t����A���Y,�2��{.\@�;e}$���3րh��\zL0� �a��sj����<k-��
��`x�^��VXI��.�4%dJ��7��1۠v�ڃFL��gCT���Vn����|Tߺn��gʚ��#�$�Ai�3˦�]����z������ܓ�Ü��3Q� J���A�m��4�����ܫM��&�OjM�]*yoqVགؼ�mC8U3�T�k�53�,�:�W4�}8�����w��B����}�~᥽�~�$G�F�u��C�A��Ӑ|u�?��6���y�U�k-�
"�BE�"eh⤞hS�^���q�B=�H�N 	��v��d��O�a�V\N�ˊ_D�R���TD���#	�T�P;/�K�0�����,l0r&�CK���`%�HN[��4�}wl�w�J{��� f�-�f�%}8w��왗��}>-�5m i}ë�ff$�Z�o�P��}<.ڳT����#Z20A���2�K�.�>M�%���R(u$~@x52��N�qjy�8܄���qi�f����;�	
�Q�O*���*e�����*�&RT �����o�R�� ��I0�[u�4�}f�?�����'��ino(�^RX�Φ�w&�J�$c@�5`*퀆�x������ҿ�'��:_�wp5�B�$̧�wL5�t̾{(�<�0B����}���l h���|�v7��e��!o�|a�uM=�'8
�H_~:w!��"<綾�
�!p;$zg5�c'�`[�U��y�Txy���H�gZ���ppZ����m�[]\S�{�˞��B�˖�~g	N-+q��";�Ue%��R?5�̯��$�Q�=7=����
8�5�!:Jd��\:(MMۡKL�G����-�����ݝ"!M�ߛ�E�,�S�fC�Y���v�47x��!�Fv�>sX�MU���el��s��Z�f�b�1�s��bO���{�1��]U�QvM��l�T�m߲EٝM �fjR+n}�K-O��2l�6�%��,o����<�7�J�'y�q,�]'z�mI� PA#�{�f^X����4R��J�{�A�Ɍ湚����I�q�<�ޔܣ.`A6��Q�/[�_�������Xs/
j�0!���\H͗@�y����~uiź�#��H4!e���8l�����&4���+�*�'P!d��٠��u��򠒋�M�z�:}��Q��n!���/J�W�<�����dˍqu��l0����<c�._I��'��ȑD�׳�`cP��������o�X�ʲ�� �1���jw,�X0W��FP��'ف�!lY�8��howV��Iȅ�aU.��$���ݧzЍ뇢�X��	O�NGF�)$ܢFF���=��v�YId�%Oh���k�̀��pV��`�i�I��$4^b� ;$_�$�ײ���v�}��sp&�>�C�%���k�u.vRߋ��>��v���g��t��Pb�FG��M�D^R�ڸ �YC&�Tύ]*��Z���jN(�0Q.~��8㺽��cĠ�x�.]����EC��M<Y���|���.�R�Ip�[�7ب�V��㸦��� ��p+-�
|�O��ʋ%4�t��?�pBJ�A�d�6A��0��R���gqN�$l��":���
1�Z��m�s��q���ھ+-~��qք�I�xB��9��iַ_������W;H�q�Dl��R��=����X���ot|5�#��O����q J
�C�#(��L��弊-Z~dtt���ؠB�hs�v*(6y�a�y�fh�V�s�+`Ξ��vnO_3&���������0.��H+_��>ݽ���N�ߋX�b��e�+�)Z/9[�<y?_����� �0�D�7�����t�}�w�h�M�`
[�iՔC�@p�톈>���4�,� /�@�rVQkՏǃ����&�v�[�Q�v*��`
GC��"\��V���`�H��ܑ�5�~�p��V�#���
;|�M=���ك}��Q�/LC*['RSt봅�j�e��ı���Ѯ��V�/���f�wp"��b��e?l��>��u��Kd�e���À
�u�\�<�$:朗7��[	���V3�e���b��=qk-lb��E�꫻k�mM�(b�,K��#�u�95��on���?@Q�Iu��[/�M�Yz�dY��x �MaV��8�~Xj �/x.�i�!��p��-Ur�G��t���5��"kz�M@->m�U|�J��V?�ޛ��E�G��Q����F/�O�o��)jJ	J����:�x��w8�י�[���QXt[�B�Z���ac�Qm����'���T��OQ��R��hu�t��<���ײ����)��p�)Կ���N&�w���8I��T�퉠�&SI̰�4q���ؐ�a�?�b-k��	�����&��}`6	�`�Ҷ��>+[ٓ��<�� ��b%h�b-zD�A�E�J��E�]���38���e����p@��.�J�gl��������t�P�O�N���S��wpn�<�=���T;Mb"~��q8a�H:Դ۞�o0��)�#`6�p�2q����R�5�/И�R��I�Wj}0�Ừ����1?�ku"����O�y���8��k\>�2p!t'��Q��6&	�%^l�_�/�}cv��*����MM=7� u��)�W���~�m���WC����&i@��RW6�E���$+h���1�x�����#u�"���?�R����m�u�!�G�b!����M��f)vF��Ò�9Y�"i���7�s����b�Sl@Ip!$�PGP���#GBrm${����U��r��ǉц��Z��y��(a+�w���o�
�T��]ө#	��}��r_ޮ:}�u�c��2oc�ɠt����W�!��}18�וFK<�i�P��_��[2	S�I?�����k&�+X�#fZ�1�C���Ǘ|Z���<���^���o2G"Q������� &Z��@<����� �䏈/�������qP����:%���� �t�)	%�)�~	%|T��^��0���9��϶Nt`�����HHk�:9^ĉy[�|[�> ���+�c��p,5\J�K0~�-� �?,���������{6A�%*3�O@�hEY"��-���o3�ǡ.O@��z�� *��G.Nh8���r�&8�A�[Q��@��,��[��Z���"9,��R���$�yp�J��5
2.���Obv�RFj_E��X��jP5]�}Pl�Ta�kg��x�K��4ic�|�����,۴�*�[}*����� y���]o��5�?�n��M'�M�W������s�^�>�����׭R.q��+H�q�m+��/��X��z�<Ym�F�Q�M�vTӂ��d#�s�H��`~�ejdjWh�zJ�#n�D.8�d)���|W2�X���N�����|���e� ���G�.ԋiؘO�s�����>��_�,��s ��XZ�n	��9~���t|�y^�_.�k���]�r�P)`z���C�GT?��	C�|D+.FH��.��q.���B��������L��*b����ˁ����Tb�pS��^�N�
�k���:ל�t�n
t��s��Tݓc�����Ox"�]_���Rps ��5r��eFFc?��͒Ť��>[��Opڝ�	R"c���np�pMW]��t�Gj��ft�?Y�`�*ih�R�;���r��co,B� -�UL��(�Z���We�Q��͙f6���<\�f�gU��Gz�|���<�-K������l9]ښ��a�7���~B��;��4�h���w�ƱP�
aU{�5�8���Xș�|�j�hۀh<�FI^��J�����.���C��Z�}��^�	v@�(�j���|Q|����Q/�ذGqU�B�"@�'����0L+�����L#!�&���7C�I��.�V�6��]5��9&��ay�.l�+9���_D+Sj���､8xX
9Ś;�� @��#l*g�U��-F�Y��8e��M��^{��Px3pI���}�kqa���ׅ�VA��psF҉�kk�v���(�7���x�2�=,@ҿ̔a)������x����.��yq�{�
��Sm����n��Ù��*����1/A4D�ў������ZD,j�ZMW���h ���S�ɥ��`������S�`md+ "+�oDL�l"����2K]������YU�zB.�3s��5�`V6�X���#�I�pv:U��G��`��`?��" �~���^�,�%�^?+OWȾ�?ñ'�U�Y-�p�^�L)�o��(iX	�3f�M37p�m��~�Ƈ�����Z��,:5�oc�	���3�"���F٭,�z5h�02;�T0��a�dv�~�#���n��!W��w��c���y��"�C܉��G��c�YUp]<k=��Fl$�t�2K����pp�R���xj���Ka��>W�	������� �⌄R�}����-������5V��`^�j�m ��ꆸqJ������y�]]�5���6@ׁ\� L����<(�$���l)���&�q�hiRoO#�i�8v���׌�	�H�]����&�4�h?�b�|v}Ү'���4�N"�����f�5�#�oa�;��O/<��!n�%�g�����,�=����� w�6&&����e	ha׫����)�xc&{ؑ�D��ߔaؽ|h���j9��x�������N)e�@J� a%�� � ^�]+2���Et~Z�����9n,���bTL$>:�)���4"���.���Y;����C#���xp{A��?���LA1f�Nnq]��~���,}W`
�m�{���5�ˊN���ajH�R*��
��h��N���3�9�.ʄ�sZN��X�RE��`���R��V } Щ��={��ӛ>;L�)-���*�aea+�r�C�x��F��Е�PL��4T���H�rT��r6�҇yB�`��+�7�b��s�vf+�Jl>���@�$&���k���/|8�G�{� X �"=tE�X�,����_=����*p�m2������0'�YU�EoN��=D?�m�!m�/&���'��8�B���sٟAP�Ӊ�VK�>�w'E���@��H�;V�5#a��,��,��a*i]���Cd����`�U}N:Fr��X��i�wo��}=�O�0�Cw�� ��?����`�r�1�M(����5h�df�nʹ.���	��qUA}��CL��6x���Y嗺+��k�Ky9�!�p�A@o*�Gϸ����l\NQi��:�����G�o������29oB�%�h���R�w,Ta��-aa*tl+��ﲼ٨��#&��W����c��|J>��ǵ�3��6KE�XZk�=���������jJ�a�Z굆R��K)$�+b�@E����'�m����۬/6����ni1�W��)�^q}�%���gb]?��y=�fb>��������nCB߳������wK�C)6�g%WU;�UX��h�½�S+�99�]�>�x����O�n�?,�î�F��(1���:��v��5Y�ò~Y����V�UM�o��Ao�4x�8/#*0:��c2ڏ����0�M��"?
r$b�}�5-e������7�V���m�0��nl>ٝ��t�*�Xi�&�ɢr^�<ZS�n!c�0Ewi��Ws�����>���T*>O�Zw���#��)�Ε(���'Ux#��[��m�7ͦ�lQ��Z��e�m��o8�F���Y�"�K���:ZZ0��;���f��.��be���Y`�KY"���;�o?�}����ͪ�	���(Ջ�	����'����i�:�����Y�:q@�.'@���3�JKsOh�����
͕^}ѫ�P>τ�d�ƣLs�-��-p��ǻ�Kx#┆�p�}��zk���fC��$��ﱵv|u=-]��<l�D�߃-s�S���b�S;�P68��vߌ��(դ��������q�,N'F�[ur&K�s
*��cBn�7�g��E.��T{�J#���R����A��E�k�~����+ۊ)�
Ar ܠ��b���&�3Sj�K_`/�P��s�Ls|X���~,��d�*�7�BX�bi��&ƿ�*�Ρ?0�}\3�6q�=������V��b������5���I>���� �nzX��!"� �M���(�R�>(Ў���d �B����)_�#�O�/����E��:����ϝ97A(�W���Y�G5�l���A�齢5�酥s*-�����u�t+�16�p��v������D�nN ��+^��Lf_4�~ ���Rb䍕�iKy]УX�ĺ~�b@�iZ����۠�������w�Qb�������%_�J,�]�8.j���'#���Nt��"o�W�p��k^6�
l��B�Q���7q�/ �
`P!��@�9i��y��;t�0�I�l:����1n�ӥ�4 ��S���iP�]}^l���6%��˃o���ꥶ�B��$B�M�;�/�e0�>u\�K���`0�u�s"уf����	-��9cW-����׺�^u�A�trlQ(C%�R+��f3���F埬1����.9}|&=Oڑ;���XU�5^3u��G�����7@�a�2�U��,�u�GL��O��pA�!h��Yb�t�z}L�i/�q͹�uN��}��b���A�Ez7 �j�0������ x�;�ɛ���ܝf���)�*�G'�<��K��K&zZ�Ӭ4o�s����g�;��f�)k|���2�o.�ٖ��&<A�i=���?����~(��]UB����>F"��[T�}1�\P=zd:���G�Ü^���`GSVk���$��x�"zx�~ܒ�&�]Yu>�a�)��I�{]�)_� ��f�Ĝj��S���n�D��fʩj||i�mF�Քߜ��$&틫��8��lۖ*�P_�X|x��3O���Iܺ�h�Ʀ�yW��Ӵ�qӮ�<
���]m��΄�v橢���ś>�c<N�>+Y}K��E`��>���ϥ���1��I� �"̑m\�u���5L��"�[��+�Q�#�������6^�3eX��޷:�~w�
���J(<0�7{���l�"�u��8N�l:w�)�#�Y;����D^n��-	�P&��4l���b�-]�N��M�^Ge��~R���*eJ�`c���5�j�R.�+�����4x}r �]z����[QdL��/o���bL�`f}%nT.�&'�+��~���P��J����}��L�!�7k��7�s��3}��MT�P�
��Xˤ��/��{����÷���h|��SwO�V�lV�XyL$eƺ���ض$%���6���g;��ǀ"fpJ�ѢM�|�Ȑ@�,"��͒}��]+����6��`��V��V���7�Wc�t��_��.t64��Z�"�%���~�3�`�=�,
�;�^�[�~��`��Up�l�ht�i3*%�3�,��x�=F���fR�?%���
����"����+*S��E��S',�՘�����2����l@���0)��'��>���w�Y4�/e�LdA�$�4�sr���	�*�f��������o�-ɮ�����.���������$��-��%��!�-s�>�	�8X�=���n,��X���;��m?[W{'��cK���yqZę�=_te�A����8���ѿ|v� ��5�:�wB��;��﫽>�ц����~O���Du�B�J�j�%�6�7��^-?�b�l�T~ ��O��P}[%#C�]�O��X�P��,��^
l����T��HY!�H���?|`�6h����tG��Y��r_M�}�*�*�̾tW�C���4��n��,��-9�0Z"bD������'�ю.���(,jX���M�~[���a��Y(z)"3%I� 9��vql��ӛ��P��ڇuV���]�auё�,��ڪ@��|��y�wQ{��|��;����8���H�s^eI�J�����^�%3 ˙#��=1ݚ3���2s�����<�e�TS�
M��fKY\n�M�X���0&wV2R��@p��3�XG�4���ڹ+n�ז�IF9�HE`��f�|����L%��z���b���G�^�|�*8~gI>4�`r�s.�yc�ԯ�W��!�I��Ut����u�L�Wc�%djx�5����$��Z��E-�6��#_�ȧ)�)[wXh�.m�x�ۦ��*�9ڻ��bϳ"l��Ã��ިCȀ����{�x_� �'-C�����p�wL]����4���`K�*��޴���RoIGl����q*��@|�	\�,�#�0���"��	���}O�d���6u��]R9�a���̕��eI��>=F�8�K�;Ȋ-� ��?��o�3���>��Uw�y�#�0���R&�6����·I�I��Xhݨ%���/�p�N+��b�y�bs͆W�&�%���HS�݌	���!�!^~3��k'���o��nT-�(Ҙ%������Q@�ݾf���P�؎N�	����'X�I���w�O�O����>Dj��
�+8�-��
{F��a��Y(�H����}�$�,m5���)��L^o/@�ݿ�4�2��R�7[��yH�z�����c2a��S��� Df��V:[�v���d8ʚ��gE�D7