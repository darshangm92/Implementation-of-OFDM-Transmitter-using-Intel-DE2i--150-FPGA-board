��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����;镬���IӒ��wf�����`��ONl�C��>�u�0�w�S.Th�dMy�|�����i?���$��	n#��͈���jUl�f�4�lR�x��6r��X��SH��l�Md��v��L�����<e�"��!��%���xv4Ü�<��m �ڰ,�f<������BE/r}mq�`bӷ1L�F$F��+m����Փ\��N/:8�'g���_�K\ϥ�
7�J��Cv�4��!��bcL;V����94���6�c�I�0�v!{:�z|���t��~�Y^�E���r^�#�&d�
D��1+7y��ϳS�j�_��3���y�z#��%p8�����2b��!�1�%��8mE�y�v���Px_�%Cȑ����K��H�Xxt6r�|L�c'��sۆ��F{59U�ɼ�n&	��-ѕ(�d��OAa��@3�����܆ϋ�)K*wa׊g�9AM��`��U��s:k-Mn�K
1���PW�9�L�H	�W�!l���"c)�"ھ1���VZR�3ׇ��rU���hFBj?�+Z�qL8�-\���?�@Gfl�
�2A�4�o�nM` y��ݿ w��D݇ TƜ�h��r^���>�'
�2��S+�2{?�����`�V�HeY!�� �i���xj���7�g���ഊ=��u���=htW���D��=�N]�$iCN�OFE���=�6��-B��o�G)*վ�|�sg���E
:�dVY�b����-ځ�Èj��Ke2�]�uhfU��.¢x]4$r�귪
�G~�UB��P!�ګ�C��g�y�����ϫ�\�i���-Wc1K�z�\6�G�^���D֥�:rbNEg�������wl�]�~�ד_��>`��O0���S�q�����]��c_��Kn�dd=L�G��Se��^�%�2�l�N(���D����Ja�{@�0E���r���,����ˊ���4���r���_�<1�Ss|��Y�W� Q6RM��� ��w�����zA�G�P���c.�( ���!�$�T��𖮒V!��"�~a˵O:F�W5�0�Y�v�۱�\��G.��S?GH���^(�@R����S����pj�j�i��P�1]*��z�Q��J�x��ck��`��6����G:|��#�j}��E���z�=�)cӘ�A,�� �e�%����~W�br�M*��/��\J5L��+O���'U�Q�[H!0�j�'�Is�����ײ�q��ʏ�� ��*Գ�)�d��Z �EAګ�UN�y��I�X�Ќ(�ܬ�Gm���~Q��f�{�R_��8��64?�Һ˛;k�`%4� Z�jOl5a�M�.['D��R�ڤܳ� }����{c�<�p/@�)�!���C� 6=�d�y�{G8�|����L��>�Z��h��m4'ʅr��"��MQ�3<Z [p}ma�oh����ȕ�E'#������T��%�����*��g� �R)����jҏr��|�r��Q~䟘�7�{b&D5Z��j����6�?�)K���y5y�?� :X��VK�c��R��Ձ޴z�xQ��3��[�����w0�rE΄�m�:�O�6��ϯ��]�d9�h5Y�e�����\�L��B��mk�!c�nq��4	׻FB�㸄�$�����t�1���/��1��:"����N&��� ��9+�Ѓ;a����t	L�H��M��d�Q]m3���LVb�i�	C^W���8�(*VTC!�$`�@�0����bN�NG� K�K����d&���]x�T����0|s���x��P��1��T�g�ad����@T8�#X���N�&�?E_�Q�d�E#��Cr��1qyF^�34	K�br*�W�WN � �DR<�0�7�A
TO���ȓ�{k�y%��c��9_�ע��?M��[}�)�ب��IKv$~�R��c��,b3�������� ��n�HT7sA�����S�]�W�ؓ=`�ꭶ
��y�t'�f>y����2��Ѣ�^�W�G���L��Zֲ���nt	ګ�����Wή���I�쵅/�G�V��>�
-�b����s� 5�5�3��{I+�`n�c@ ��8��W8�W*�k+э������
@���?��:
h��I�:c<B=�\�P[��7y�rQxI�q�r9˝�I����fͽky��J1��
es��-��*`��e��W�a#5�pKu�F� ��|�̛��11^Fs�P��3O�h�p1iTsh�������^��p��NI�S�������{�s
 ڸ$8��)>d��*�fG�X�2>w�E��[e\
��̅c�.�����i���8��x�
�l�� Z\`�ඡIA&�ʮ��drS�xd�"���z+��̼�S�}fy\/�̏�
��Z�z�4S�.���_��B1I�nV�p�P���҆M�X������,�eq�b1�#������,Y~��qA���X����8Su��P�!k����F_�T>\3��!dɍ!�os���1�y��-++WP�s_���%�G�$�}��4��+�P�d�ؤ�������}��!$|
R$]�E�U
����8�^eI�3 ���WiA���@���s@�^PB.���V�����q��^��a��#l�0%����%�;{ዩ���R�V#�m�)��*��s$�\��!uP:���z��'6�,� F�mW�D;70	D���i�.*��7�O�']�]���@W�*�ԆD͘碉��rE��Ǩ���
}��Hٌw�=�i��7��Ӱ�#8X�$�,�Hr�+D��I��]|��<��9v~vB(�Gy��v91�O�7���TB8f1ؙ���A1^��F�dlW���O�"��"��he�A������(��2<J8�3O�V�]ە�=�
Y�]�4�������c�*�E<�m&�<]o��_	�O��F6 �GH\��l��4�8��9�0�F"��f�ہ:J�ߚ�Y�ҍ���S�R���>�L׺��?D~�t'��?�(��Z�*��u����1�j�!�t��,(�x^d���x�lhI]sAn#y��d��e#����#e0��H�˂&��]������t��81�Ʒ�\���DG˅�����\c�n`��޺�c��h�X«8)�\��"���'��X�&_�6)������h@ֲ���8A;����A�mT�`��y;l�//M�<�:dsڣ7�{��G���C��e{+Bъ��qm���x���U7��H�l���0�8�����4�%�S�1Ń�\����H�&����1mtsc�}˧�D���1��|�[�;���-�c�d�/�ϊh��k�g��Iu�̶���4/�tH8�����`k~(H�1�z��	KϠ�\n��p�L,K�G��%��g��D����� &YD"�l8�2R&��5��|�z0�}G8��N�]Ă����W�)�W�ư���Cd�8B���}yo�0� ���FH��������2�����<x�;�H��y�Sl�.�&h 1��5<����h�d��-�h�v�����}�3�M�T��#�v3�2�0���Ȁ5EG�$٢w@I�r�/Mw��	i���%L6���n��ӏe<0&_����7{�r��X�P��l�_Σ���"��5J�ޞ��<B�z�(B��-�!�l�IiF+�-��J��d"e���*�"ZZ.���J��I:�
�	�a	@�"߆����0}�L�����m]�K<:�a`"gk|l���D�6>:-y29�2n�ڃFӓd��"���*��[����O�z�V$K���8N������4�m�9� �C��f�he��H8��sLN;��,]�Jx>��'�\�|�w9*��*R�n��#=�tw��6?v� v�)�}`Mn��� ��Y24}�V�2>|g)};��d$��(87�����׭w��^z��v���$RCXh���g�t�'J@� �Wq)��j��l��q?�_{$��X�Q������d��j�}:�A˔��/,Dl�b�L}u�5(��F���s��,o2 6�4����D��?������Eg
ʯ�����6>�x���<N��A/wG�	 :�1���l�;�(�Ŵ���>x�Pa;�	�Կ!\��/��Dov��Ϙ�A6��NP��_�hU`��u�E��2�%U���<��H��F���#@�ID1�f��r	�IGM��u"_,tH̎f�X!��|��j�_e��!���:�c�d!��Fh��/����\�?�O}M��}�G�ǡ	��s�2�$��8��UauӔ`�أ��������r��#�~ډ����
P}�Y;
�N1g�þ�17�(�=�%�:�[,�>��pj�*>t��{}W��@Ms.-�{2�醶��'�Es�Bl�^r�����k1\%ti����0Hv����i}>h��f]��-�v2���X�' �$6���e�Ұ@��9�6q�4M�K����D��
���;N�������Str�m�l�D����!��!��ɄK]���\�)���cL r�`n�>@Ҙ��ʌ���&i�6�V�����Yk�M�6��qf�ט _�hR��؄w2�'ׅ!�{���d�#%)���3*��C����C�撅Ve��U��M�2����8}^��sr��npXn!o��v�����<B��3����`en�|s�1;	Ѭ
�jV,N����R���_�:`�y�a/��=bZXF��Qo�l��!·c��_M�d$4upl�ܸ_Jq�����u|W�M;�s���i���&����yZ�,;3�AG���U����xe}��&)�9s�=)���Bn؅�m��[��zIMe��`���-Tǳz�M���J���N�
I_Yp����K uW�l2�Q�nĽ�\���'��R[t�X⵿���R�@Y�J{�FQ^�q��u���W2�]�6Q�)sX�"�{y��H�$������,�"E�-��O%	7���wWt��2�-�"�e�bӕҵ��I��V�@MI�D�S������ÔEж�Px{$���t�H}�c���-����1�&0m�z�r�3�7˃�Yg>9,�$Q^0�����Z1�fU�<#�L�c�<��Kl���i��'S��""ч�ڔ'��	k0m��re>ʣO?F�/��(��5P�YX0ν%��R���K7�4Nqc��Z�c����峴��rT��D��zA)w�5Ȗq`/�7G�]��!�:(z��4�J���Ym�j���Y�8~�2�	p�E�x��bo�%��%H�.���Q��_�Nlݶ�t���r/p�E`�[ܤ�,��*����7��bđ�zXs�'�A����t�!��6&'�]�a_\`̩h�Y&.�͓��`{)�,:�7g}���@���l�r��uwGR�a���N��G��R����Ă���t�q|;��za�C'/@�7):��v�[]��8�O����t��u1�E���9Ѿ`�bVm���~l��&BTȨ�*6�FG���O�%ǣ���_A;���8��NM��ۛ׻lS�V�,~����2E{���u%�8`���:2���9��H̥)��F��s����4^��z��<.�f19?BR���2�Y���wA�?y��G��d��y����M��%����m�vt�aDpU
3�8:}��d"Rݎ3�y�� ��Hh��"7��'���3O;���5��d�L����LNr�kEPW�������;}�pSo�G�iEh�sH2�n�U�p[j�z����H�K��G�g�	EkS�!>��Q���W�^��E�[�^{�<8S-�ɻ�A��%XT)g������>"	}��w%�{jq|������a�3�2�P8����Y{�f'��\��+�R6��O>�����^ c怫�PCE�=I�}�࿘w��^�(���ߧԋ��H���' @)\#��0����g;n-ݨG����aV�_	��������X'lodZv�I�_x\?4��4�o��H��ZRO��_l��vf��� ����|j�j���+&n _f8�h+;EM�C���{�m�/���I?;׀?I:*�-%�u�?�^}/���8c�-����"⏰*�{4:�e,Ͷ�>�b� ��X����hd��뿲���WMy�7oD`B��b��#�.��%����:'u}��*�U8�ģB*��F(�|rp^Ё<߈��`���%�ޓ�7̨P��G�����h��e0w\����]׶��
�M��fq,~��~}�q�
��Fu�j�c��VhH�j���w�ifC�u���1,�|����H�����=�=+�+�#�]B�$�>z�}G�>��.
�f+V���'�U'�$хc�]�~��t����`}����´�J�MOj,���ʣJ���e'+�	��VC�I����5ǆ�ަa[x�R�������" M3�������>��D����=���	(Â�e�Eɷ44ϼ^Aڣ����n���(	R\oj
Q�gl<J�� \r[Gu���'nU��xɍ�G~�qIG?�W�9ྈ6��B�M�l/��"�������}��'4�a�+s�~����y�����.���w=p�I�3��i���5�E6w沸+H����G��3��Nd�RT�S�U�1s[У�M�.�r:�I�$4�wn�%A���!;�?�dp�hP�[Gx�##P�ތo�~�1��l_��Vym�}t�5�����r���ΩͰ���C��E��z/(�F�ޑ�~A���E# � }3#�)a.:�Bt��������C����X�/�*�n��<ix=�p���k�#m�[5�J�)��h+��?(�l-�(}���
� �	|[,�I��a��o[��:y͛"�0�cU�.����O�=0����(�l���?�%��X�)�]�A�}bsN��ن�b���
��ʸ�6׸n$��E��4 ��W c��>0�>�����~�S�,q0J�la�3?Y��9f�{!���Z�<�9>q��0�Ϊjf�J���2�JZfo��x5
��lm;�r^	�h��<�㪿}+�JK#XX0�~�IID�GLT��`"�Ä��� �H�c�W�qʛ�q�ee}��9jsd���9'�s��������� aN�Ӿ,���%��G9�WّC�G��)b5�)]!�8:w� �^>���:��D�SQ�["�s�������m�n�W�ń�����,Cp���F[+�;cI٭�������Ð>��i����I-�l唵����Gk��f.�It�Z�?�m��=-��j�`���y�+���N���EV�!�Rpն��AЭ�e��?����Y�P/�❤m���T�:;��-�i:�~j��6ŘdY P3�{�<��TDa�Hxz�F�2�#vw����0��>��y?�����!�\\Ȕ7e�Ѿ1�����t#��|�� 7ғZ�oa̢iC1��|PY��?K������xc�"�+��H�,8���9���ِ�F��|�y���:U�b���8��~��ơV�J����e���(�(��n����������Cm��K럐�B�L�9�_a�9���w-K���	6R9C�PY�5f��o�.m�.Y�i��H@J�{@_�r��y��O-�8`��q��H�k��v��j�����'���[��K���{�F<��:�l��`�f2�#kj=s�W�N���<U�(���}w܆ئe���g�!E6�SF�1]�Q_��Ę(����ϊ�JPJ��4�����:�2�iG(41���]M΂TC��:)5��bVk�m�*HG������� ����˗�K��,;�}2m�r��u��6��O�)��<q�S���aQBԁ�(�#�����.C�T[��j�S�Sk�4�u���%�G��P��!O �D���&^)���H#�|�&[� �@�伎�&`��"�;�i<����O�j!��=�vwwb0���R�>g|�ִ��=:��#���;��B�����I_��h1pNP1GT��A/����jk�Rai4����a�x��ik��זN��?��C�����O���=R4=�XI*�-�4:�z�%4`�����3�5��y^�ڞ��GF%���
C��]�&�����Ȃ��O�����v#��СI׶�E|"��&���f&�����������ߋA29�YS�ՌM���A��S�
������n��U[}t�w=VQ�α��#�0�4%�i�w�v�l'�6vVR��`l�Bu�Wx@w"���H�|<u�ȳ|�}����h	����]��is�)�C�sTY�����V����.h��#R��?�y��6����Z!�U�ص��G�A�\��Z�&�k:�=^�Ғ3]c{u�aa�s�n���3���T$��]6C��`p����u7�M��#=�ە'
�x�q_��+8�ؾ���l��gd�Tq��E�,gR@}N��/wL��p���龕��� ���1@P��ϥ�W���1���:����,���ٵہ:�6�� ��hVӜ�W��49�t8���bS�����	����C�Ǽ
�KH6��=ݦn�Hi�z��8,����֘����ŵ��lmm��>�\��y�T'ز$���zQT֫�@]�eaq�fE n��eVC3��z��m��$`_OY}V�6���8YU9<}#�רJ� B�ҙ_e�R��CB^��s�<l�7����QF����R�x4��`N7I�� Ze�0��
��&\�(��I�Rd�8�F��fW�������kk@JkF$�� ���-c����*s�f������7�PƜ*�Pg'�ȭ�A�x5T8�@�ꎻ$%��M<,���Vp��a����ڿ_F}�zG����7�[+�����ݘc~kz��:~v�����-mPC1�j�hwe��7ȏ�M�&M^��R$h0~Ԋ@,*C�j�7G�ףQ�.�sgΆ��N�qC�d=��)g.�K���/c����,y��/3^�5�E:���|�XH���|��@�b�k��)KbA|�P���P����g=�R:x�l�t��s��T�l�V���������'>B��	�f�"��6�m4���"�́W�I�L�0�����d�Ij������<	��p�s��S?9kA_~�v�t�Ot����΁�dk6e30w�&�^�Φ��'m�k'n87W�}��Z�ap�nx.�.<�#��Dc�ͪ���\g��K���&X���\���{�y^��FV�:�k��;|;$�8OHV]HW��K�9Y\����Y8p�Xc��Ѐ
��'m��&�k��[��bz�Ҡ#�l>�E�?1�o�g1
��[�f���`��/=�7F&CP�����'+5�b7����0����R����?&_�z,�_�� ��핁ޕ3��u u""Ӳ�S�W���Z	-�v�D,U�����a�U�!]��k��_��u��R'@n��+S�UZ�D��=��g|k}>_[E�G�ʤN~��z����� �Ϲc����&(���992�W�<�Y�Ł,��8�'�#�5�+Ϣ�	����U<K���Dn�V�_�pqC�0���5[�}��`��}޿�e��h����������I\�w���g>��V"����Fa�X��}1,~Q.w�!NBi- ����� �xΏsW���k�G�qj���B�j��JS!t��z�hO�6km�p���Ke�a���/wz5�z_&������ˆ�����ò�x���e�����	�51ت��i��Ɠ��CN��sǡ���s@���[T��Gя�5_���E��a��ld��@�H�����,��� у�b_�1$�>I�'d{������?�	x���ge:JՔ�*������Ć�|���o*#���C�8�h.Ϟ$����?��R�:X4 �Jr����@<s��n ���Vt������
uM8a�/���@�	u�C����!��?y@t�=~x�0�O��Zd{a�S|��=N��R����tP��d^���ƻ$�ɌW!�������w����N�^~�B�&q����d�����-�����eIU:��/�~����_{ף����(h[� %��<�P�*+�������[�����9��"ƪ��~L���e�M#
���V��ۘ*�+�� �M�P���p^���fST��1��t$�9��m� ��xj�'Z΂<,!w���ÆD�1�ZK�c��̲!$/Q��K�r ��a/�_��e������i����̈́��LS��y)_�U�Ek����<�z)1Q��J�z��)����l� �` ��?:;�5�����&5����'���qe�z��s)-�5�U�!͂W[����' �\����%U,j1VK��X{dA��C���8�P4�
�z|�_�b4�Q�zH�8��u ��|�>**�Bn���|~�U�:[H��s��������i��� ��y�홝^C��1f�Ys:,N�? ^R�y����5�g�����~�����w��|��=��9B�3��`lu[���R/S%#�ӣYxt԰���ҕ�!�מO��J`�m<�3Q�a2�L�[<];M>	�^W��$؂'	H]���1���l^��2��ˣ�6)x�s�ەt��,�Ƨg��Q؁�J��s��T�}�n�J�7�=����=��I�VT!ē��s0u�~�мL���F��})Q��Yv$:����g(H:h���.�B�`J�iry+Ǳ+��� �L�]�*�E��Q�S���*%�K	MF!`l��@6(g�k�
 �_U����tFͳ��B�0�`���V�k!�n7z�9Ri �I����r��*��*[����今YN�W#��N�gھ�.��v�5�1q��8+~�**�f%͖(�UP��9kBp��:�`�z=ֺ�i���h1�d(�B:�D �GEշ|Y�'��f �e��鞘T�����C��C3���pY��d>�or�!N�b��X	��)n��p��R^(7]k�7����1�b�u,AUX�O�.�F[��u��1rR��7r��銰FY��;�D&'gGT�PQV��P�ݿE�y��>�p���/D���0��y5D�O*0}��k��9����3��W����Д�����ٴ��gvv"�PҚ�J�����	,�kB�7�M��z�q����hz�@��!g4_>�܈�bH~q/�y��YJ��T�&���8��㡈aX1mӄ �9����������V�Za��e���M����#t��NM��kbg�l�/R�So�I�D�j�XIc���T������R��Ѐ�h��J�"'�N�B�WX0��a�x� ��?D/\�!�{s�,�L�h��'TK{�}�<B��f�8`�'`��7�4��b����ץA��W�BA��|��&dpc�L�G��1؅��g*�A��)n�nK��&�_"[�z"�=:���,�a�]�4��<qQi��D��4��	�ĵ�bZ�x1<��FW^�JM[^�wơT�-�g���u���I>���8I"YP�l�E�
8����'��{%Mk�u�7l(L������F�?���s<�ۉ����~y�w0�nh�Dj؉�9��ޔ�C�fZ	g`QϤ�{�E�E;�?i��pL�I[�_����i��t��B_y3t}��~и��i]�[��g���gI�i���%����Fz.Luү��f�8mF�3K���~mWH����L�25��}ԛ�������$���K�E����"t$��́o X��L!��;�K�á.�Pl�~?�FU���ٜd�{���_{oY6� F`��e�M�� 0�o�.�|�R�93T������������^�>(B_�4no�a/�*�+��]��o�{W�P�*SN$[6̭-�6�����^P���N��m��~�����?��\U
���)�榷��J��Y��[$!��-\�W��6��A�M�M*o;x�T��m�v��'i�=���p� �ۦ�.l�m>KJ��۩q��� ��slo�PbR7f�<H.T�~+(�2�Th�9E�+��ʑWh��`��۫r�3W|P�����afu[�AV�V^���eVU�yc����/]^e�=-ڥO��!��,&�G���8]�������);fMI����g����ܪL�dcҌ��h0J���ƬwF1��ԴbK�泞r����S����hEs�9�9�@�!�݋����54���O�9�\�_���V�� Rq0?"!�m��/�_muza�օ�\+�ƥJ���Q<�3�V�_vҚ�>IcVA�F��8a+�~i�o����S���}l|�L)�>T~��#���"����Ql�	j�����64=n<6c�b�a�be|�r�Bju������+r��6!ꄑ�\�v;ՃA$�Q���L�g4���콐2v����["��]N��Ha�ΪLu������5�(C�������RN>����\�MI6uFd�q�&�~&3.��j
��%��a�񤄝��o�`�����;d�^�敼י�qZ�6�J�]�P�Iᣥ
e����m�>�ٷ2R�_�\�kW�����\�B���yy�@ p��aL�J�)�i�� ʈ����R�Ǜ�_�dV��>�u �p��5�P=��>�c�M�����wK��i�����=�L�Y��{;�Q�$��R����.��Z*�˶�~�жB�3�;!��|��fZ���-[0�M%���ЏY���{�n��c�%�Jt�"'n�hM]j��J|.���%� ��0e��*�2Rph�P��v@K�,F�5=u�A��(�nUSփ����H��4]D���<�-l�D+�h���/�8�k�}��ή��Sqjd��-ok'K@���ݾ�I1D�N&�0*@�WC>�f�q�^�oנvK��J�L%k�z�RF�Ot9d\�k�6�SG��m���HៗEX��Mkaз�=�x���`L�ȣ�| ��.֋�"���R[�.A����V���C�R�&*�����!`�Y(�G�Q؍c�c��|kq�/���=uN��9)����FN����U+cb������¸+�Yq1�|Y�nH�a>f���[H���3�����t$b=+;�A�F� �c�R[�1�B#d0��ck�-s���7�+ȗ�W���Y���=5��k���Ib�n.��\��_��C��KCX _׏����qAs��L_v����bR����ZQ��U�-ok�N�x�%Q�����@�5��~�{�#WO(ΒRC������:�I�=A��䉀���I�U
�֯jE�,T�Z_�G ������T�hl P� d�j�W_mf���B����9���x��UL�B���"�;W�3���ۇ�:�ī��Oi>v��Re~ڭU�?�A	��ΑL�G����N��H˅"���*�ۯID$�^���M�6D��� �TSE�#�ڤ�3L�� ��a����ILy](9n}g:`Go*#�P]��y��	dHM�.�� �yp[�[n��ÿ�,!V�� υ��od��t�oО��p��`�/�[1�7�(.;9��y�ǲl�<�n�����dՏ�m�u�ˢł ١���[��/�J����!y�� v�KP�,�C���i��+�(��k����:�g�>�qˍ�e���N<5��:zu=Z}g��y����ǣ��0j�`����<���}Z(�v��[��ãD-ިAM�s����C��8@���"Á		����Vm���?�&!������7����S�X].�r��H���AϢ��6K:��U�1�L�c��<ת,b�R&n�C,Ξ���%Ir<px��g%��r�L����#���
��~-" ��B&1��Q�o�M���?ӹ�d��n���8��K4�ue�L'�|��A�߃�O>�����g��z�䕷uH}�K-,���Z��R��,���R �����!,��{[�~$���Fn���<��=�1��j?�����o�H�?{
����Qnw����g�c|��fc�Lb���ܳ�7�o�|:4<�}�<�<����j�C(���R��s�^!l<���ID|�^EMޕ7l��?Y�~��
TcM�a����\��/j�B��O%Iutr��IF��aS��F���Ԝ�u[1�[Eş�^0;��_Z�jm8?�3yֈ���B�#~�%�0]��sn.�[W�١� ŷ����>�7 ϑ@x�p�p�ѷ�>,sn�;����Y%̛��i0Lwّ45�Лw�ܣ�T0�a�҃&@"��4A��+6����L���X��>U^.�M%��B�m�x/f��|H� ��xS*:�ȕPX�����_;*��R�依��`\��[�;ko/W0�����?W5�nv:�����Вbʝ��xu��p��~��Lu���u��ՙ����C\�`z3�f5��b�6{q��NJ�`h�|���2����3���W��]ٮ�\9�r�FDS�d��RG��oCi�V0�#�g~?��V��7�tK��~FiO3B��2}њ�
���T_�E����$�l�o�O�Kt-*�"÷����?�}�x��S��y�:�Z�����R�9���Ӎ�	��vs�.2�<�҅*=DCc���(l����ꜿ�����x�2������O��F��!x����+j�vVE��2�£ɛ�˞����vE��I.|�o�ձ��^����LE�Q7Z�{�}�iP�)��V���N̥i�/Y����F'Ah��="�f6�U