��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� C|�����B�:u)=�y��P�~#�U�[�!��s�5�r�1��SaG6$��9˙��[�����͝~�	S[�\�1
�K���� )�i�D;�B�O,��0Ad��OH��uN/UX�')&(%�-����4u%g���M�D��e��t���e���������^�E��F7������Ei=�K�ӍzI�HC]��5��ńs��%8�N���c��IV�l���-P
|�o8��R&�"�4���ڸ�r����t��8*�y�
��&oi�W�^��7x�߶��]^�d�P:�϶�$iTp�%��S��XN�" ��X��MH"�y��ř{�dTF�k#�fӡ��'���Y��'L���Xm��dN�.h*�/�\!,u����bQ�y��ȃU��Aώ�Q��������ڐ@�M%	�@x�9$�v1��	��
�
`�p�$M���Ѥ��@�_*N�Z~"�Ζ�6ܾ~�8 �\�[�\�IO\�YZD�j SK+8�({b"'�~a��y">���x�S�Q=���I �I�t��"@��R�@���� 'V1YK�^�� ����NhL�oG/R�L�]$rϻ8z��o��c6�<r����L���S�vI��>�I��2�^)��#��|�t��w+�ՀmJ1����D�c,= ���uXވ��k5�����8󤥚װ��_�W�L>�l����b�"�S��a�e�����@?�����Ĺفa�i�6O��T�h�u�V�1D-+]���W`9M\�J���W,g�hm�sb���cwddފq� ̲|f�4�0Ȓ@/-3WT�K�x��᯽K��V���2n���%4!X��R T�a��!�bH׎�l���Aԕ�Fgؙ�)^�x�8����՟_��'+������d�v{�C�lCi>��C0I8zqc���[ȩ�E1U4����W�o!N0�[�̹]��7�ݚ�3�#&��#�<�����-�l�dD�i�Ս���yws�tu��e��A��!Z��7'j^�,� Q	r�ջ���*]�D�<q ���m��$<�ܚnf��Xj����&#1�K��@�1�S�ϝ��J$�36�)��f�3/�%�QS�G۫"�r�R��1U�Rh_{U�`.�>0�a����N!')�h��DX���/� �h-�&�`�Fv����^CDI)X�n�n��9��#T\-��J�rm��1���m��ܴ$ �3i�t�*�_hՄ����F ����]ʔխ��0�3'N���w��$�X��3>�,w�d�D&����TP$���-�\�2�#��i���XsA>lU�����a;����D d4�8���(8��V�x!�%.�=���hTP�����1a��[���I��f8h�ÂĻzy<�j7܉��jm���z�眛mȻETSgr�U��%r�م���(o��}v+u#���` zշq��|� �hP�����-Ƞ��>�ʤ�	�o:a\%��$��</��e��2����I)���'.[qC������8
���Yg�>��6����D1�M�' ��TӪȡ��4��� /�j�6f��4�Ȯ�y�9|q%�QW��������g�F�5|���
��;,�� )֌yTIKP�]ʽ�(�o�(��J�v��� �H8���^�� /ix�� �j����SI�.�0�x|�~n*�7A^�J��䡾�"Qi0l��M�����e�c\!3�b�W6�x��i�b������z�3�ꅃڠ �m��Yq����t��8��8�>!�e���׭.���*<�]\���L����_��G`xT��C�>\��G�vSUP(�=��� ��C�����U�V��e��+�O)@;m�w�'V�
�&a(i���q�/3�U�q�v�ߘ��q�~6��dD̹��o��(�pM��kIx�����w� T	1tمb�3����U�0����_@}�w��g.A��M�`D j��u�::�Au���5���Оݜο1����:��*|3�FB-	�A�9i�(s��]�]$�����xS��@1'�*�D��[���x�(������}�>�4vgc����߸��S�ㅨp7�]�c4ڦٯ(�>�
eS=i
�1͌D��c�Z���[_~$3����<,ٌ�4tk�n�y��"Q�m<<nw4�ʹ�x{U�N(�Qd$:�(P�r��[������ǜ�>�'���!��} ,"�;©|'�?��^\E��/�J�����[ŭS
�܀�c�8F<�n�k�v��+�U�����3i�Ū��(c�bʚdY����e�׿�&��X���r�� �FAj�Q�CLE����er����=��M�߉5<^n��S0(�Fvё�3���t�Hk�ѓI��
F�Ӊ�	6{���Ԉm�mel�"��Uc`�D:�sZ�/R	���� ��Kz��fN��; �Sx����Ļm�+�d ���.�Bq:ӓ&g��p	9(��t��G1�nK'p"��I���GJd�Z�Y=���{�1ys�߯7�/ldp,�J+<��X�k%��9Ԍ���w ����\����^t����I��<f2��!�n���\^F����'~����c�6���ɩ�����ϐ�����݈qD6Q��+��7�_��W\չ6c㵽�Wk�S������̞��"�����4;]M/�X���f���@%L�~�����{E�=��*K���s��'��L����;�@_���A�G� \�vK�P:��@މ �����pה���}s�c|�zլa�+0���|������
 ��ĄǪ
����=&{=4+>#���qz�62,h܄�w<�e+W�w�j���]�k�+�I�Nz��/�7q׃j/�%5����^�t)CDN�>ٔ���@{T��F4Q��R3I)�'��d�q�����hU�<|�N��8��O�w�A"=vS����,f\T�q�Io���Ȩ.�Aڵ�A��OK�9]P���Ӑ�?�����kgIplJ�s���W[�e��sH���Q]���伀�E3�����@r���^:���X;�l\[����N�}I�S-Bk��\^�rri�(A��D��y�*���S9N�(�h����H,n%�G��(K&U��I�k�	�-r�T��uYu惩�Z���E��U�/�7�
ro�Y$���3�m�jS]7����#�Y̟�n?�J�?��Tao��,o����atz��:�z=�:�5^��Y�puB�^E#�A��W���sΌ7&JH؜��Ozc/�)-8~����L�#�w',D�o����$ʩ����g�wD{�� [a$�J�+���E*��K>ճ�A��mD&�ex���t �M
Sv6�zz���9��_`3�)qȠ����v*���8h��^��#�4�-ŝw�~t �TV�竿���_�<jƣ�}^��:���z��\>d	i"yW���-+�sUE����n�;�[���0Ñ�Nn44r�N��5���%�W��7�O1p�V��c��Q��6ћP��a���m�[����]M>���*�|CQ�Ҁ0��J����W���Tj���8�aI��nG�}�bXT�]+fZɛ>%�\ ��z��V,�o�����#:N~�<�3��Ć����~٫LPt�J[W�=r?�V%�@�_lJ�A:��a�3�9	? �"�<4v���~�S���i���:�맥�/P�	:�$�d��͂�oEs�s/��No ��o����-
�HqC��2c�&��Ƃ	��}��a��n�S�R*�����~*�������]�#j,�`��8O��~0}����Y��F�:�*$�DS� �v�є�G�h��"ܲ�e�t�Jh[d�����y�Y�1�� �6��WHİL8���=�P��O�����옇Ggh��_֞tt�#�*|E)DfZA�����������<�d���<�6YGH�NI��'��̹�T����������d���j܊�OL�9��ԕ7�! �	7�S<f7T�BP9`�b��xH�����'����ZRy��o��y�'b�x�?��$�>�	u����Hmjo񻂹�۠6gA�8��1�]�`��������I���^.�R�#g��6	d���2��=���:�Jğ5vj���@�����!��a�]�gH>���ZbזaC��uF2���?�P!l�|�>�)vK^!�&���E��k`�C�A|,O ��7���I���c1�Gȧ�)RZ�Zmo���x�׸, y�O�j�i�6F4W֑���w�	 d�蝠��\�O���ϵ9�MA�օ��o*�Q�Xv���D'�%�(y�U�6�E[Kw:���������{
��q36�r�����5�$z"!=��=�Z|x�Z�]�G�KX�*�+��ͩ�nv��8���#z�1ӍK��P�;��9���N���%r%ձan������Պ>֮Ti�?C'�b��h�p��%q[���Q�ù�y�\侞&A'�M+(}8�AР��\EvN ̷U\��>�T�>b�/�έ�R�.��7�I���=\�rS�#W�B��J�d/ė_�d�>��ǛX�̤Û��&	��CU��8_)]�V:�B-b�G��#�n�p#S�G�\��&���������G�S-{ho�S1H�;���D̰��)&�c��.l����]�"\S}TʭT^-\Q� i�